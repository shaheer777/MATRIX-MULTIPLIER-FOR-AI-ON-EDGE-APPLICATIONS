magic
tech sky130A
magscale 1 2
timestamp 1667203070
<< obsli1 >>
rect 1104 2159 378856 477649
<< obsm1 >>
rect 14 1844 379394 477680
<< metal2 >>
rect 1306 479200 1362 480000
rect 4526 479200 4582 480000
rect 7102 479200 7158 480000
rect 9678 479200 9734 480000
rect 12254 479200 12310 480000
rect 15474 479200 15530 480000
rect 18050 479200 18106 480000
rect 20626 479200 20682 480000
rect 23846 479200 23902 480000
rect 26422 479200 26478 480000
rect 28998 479200 29054 480000
rect 31574 479200 31630 480000
rect 34794 479200 34850 480000
rect 37370 479200 37426 480000
rect 39946 479200 40002 480000
rect 42522 479200 42578 480000
rect 45742 479200 45798 480000
rect 48318 479200 48374 480000
rect 50894 479200 50950 480000
rect 53470 479200 53526 480000
rect 56690 479200 56746 480000
rect 59266 479200 59322 480000
rect 61842 479200 61898 480000
rect 65062 479200 65118 480000
rect 67638 479200 67694 480000
rect 70214 479200 70270 480000
rect 72790 479200 72846 480000
rect 76010 479200 76066 480000
rect 78586 479200 78642 480000
rect 81162 479200 81218 480000
rect 83738 479200 83794 480000
rect 86958 479200 87014 480000
rect 89534 479200 89590 480000
rect 92110 479200 92166 480000
rect 95330 479200 95386 480000
rect 97906 479200 97962 480000
rect 100482 479200 100538 480000
rect 103058 479200 103114 480000
rect 106278 479200 106334 480000
rect 108854 479200 108910 480000
rect 111430 479200 111486 480000
rect 114006 479200 114062 480000
rect 117226 479200 117282 480000
rect 119802 479200 119858 480000
rect 122378 479200 122434 480000
rect 125598 479200 125654 480000
rect 128174 479200 128230 480000
rect 130750 479200 130806 480000
rect 133326 479200 133382 480000
rect 136546 479200 136602 480000
rect 139122 479200 139178 480000
rect 141698 479200 141754 480000
rect 144274 479200 144330 480000
rect 147494 479200 147550 480000
rect 150070 479200 150126 480000
rect 152646 479200 152702 480000
rect 155222 479200 155278 480000
rect 158442 479200 158498 480000
rect 161018 479200 161074 480000
rect 163594 479200 163650 480000
rect 166814 479200 166870 480000
rect 169390 479200 169446 480000
rect 171966 479200 172022 480000
rect 174542 479200 174598 480000
rect 177762 479200 177818 480000
rect 180338 479200 180394 480000
rect 182914 479200 182970 480000
rect 185490 479200 185546 480000
rect 188710 479200 188766 480000
rect 191286 479200 191342 480000
rect 193862 479200 193918 480000
rect 197082 479200 197138 480000
rect 199658 479200 199714 480000
rect 202234 479200 202290 480000
rect 204810 479200 204866 480000
rect 208030 479200 208086 480000
rect 210606 479200 210662 480000
rect 213182 479200 213238 480000
rect 215758 479200 215814 480000
rect 218978 479200 219034 480000
rect 221554 479200 221610 480000
rect 224130 479200 224186 480000
rect 227350 479200 227406 480000
rect 229926 479200 229982 480000
rect 232502 479200 232558 480000
rect 235078 479200 235134 480000
rect 238298 479200 238354 480000
rect 240874 479200 240930 480000
rect 243450 479200 243506 480000
rect 246026 479200 246082 480000
rect 249246 479200 249302 480000
rect 251822 479200 251878 480000
rect 254398 479200 254454 480000
rect 256974 479200 257030 480000
rect 260194 479200 260250 480000
rect 262770 479200 262826 480000
rect 265346 479200 265402 480000
rect 268566 479200 268622 480000
rect 271142 479200 271198 480000
rect 273718 479200 273774 480000
rect 276294 479200 276350 480000
rect 279514 479200 279570 480000
rect 282090 479200 282146 480000
rect 284666 479200 284722 480000
rect 287242 479200 287298 480000
rect 290462 479200 290518 480000
rect 293038 479200 293094 480000
rect 295614 479200 295670 480000
rect 298834 479200 298890 480000
rect 301410 479200 301466 480000
rect 303986 479200 304042 480000
rect 306562 479200 306618 480000
rect 309782 479200 309838 480000
rect 312358 479200 312414 480000
rect 314934 479200 314990 480000
rect 317510 479200 317566 480000
rect 320730 479200 320786 480000
rect 323306 479200 323362 480000
rect 325882 479200 325938 480000
rect 329102 479200 329158 480000
rect 331678 479200 331734 480000
rect 334254 479200 334310 480000
rect 336830 479200 336886 480000
rect 340050 479200 340106 480000
rect 342626 479200 342682 480000
rect 345202 479200 345258 480000
rect 347778 479200 347834 480000
rect 350998 479200 351054 480000
rect 353574 479200 353630 480000
rect 356150 479200 356206 480000
rect 358726 479200 358782 480000
rect 361946 479200 362002 480000
rect 364522 479200 364578 480000
rect 367098 479200 367154 480000
rect 370318 479200 370374 480000
rect 372894 479200 372950 480000
rect 375470 479200 375526 480000
rect 378046 479200 378102 480000
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 7746 0 7802 800
rect 10966 0 11022 800
rect 13542 0 13598 800
rect 16118 0 16174 800
rect 18694 0 18750 800
rect 21914 0 21970 800
rect 24490 0 24546 800
rect 27066 0 27122 800
rect 29642 0 29698 800
rect 32862 0 32918 800
rect 35438 0 35494 800
rect 38014 0 38070 800
rect 41234 0 41290 800
rect 43810 0 43866 800
rect 46386 0 46442 800
rect 48962 0 49018 800
rect 52182 0 52238 800
rect 54758 0 54814 800
rect 57334 0 57390 800
rect 59910 0 59966 800
rect 63130 0 63186 800
rect 65706 0 65762 800
rect 68282 0 68338 800
rect 71502 0 71558 800
rect 74078 0 74134 800
rect 76654 0 76710 800
rect 79230 0 79286 800
rect 82450 0 82506 800
rect 85026 0 85082 800
rect 87602 0 87658 800
rect 90178 0 90234 800
rect 93398 0 93454 800
rect 95974 0 96030 800
rect 98550 0 98606 800
rect 101126 0 101182 800
rect 104346 0 104402 800
rect 106922 0 106978 800
rect 109498 0 109554 800
rect 112718 0 112774 800
rect 115294 0 115350 800
rect 117870 0 117926 800
rect 120446 0 120502 800
rect 123666 0 123722 800
rect 126242 0 126298 800
rect 128818 0 128874 800
rect 131394 0 131450 800
rect 134614 0 134670 800
rect 137190 0 137246 800
rect 139766 0 139822 800
rect 142986 0 143042 800
rect 145562 0 145618 800
rect 148138 0 148194 800
rect 150714 0 150770 800
rect 153934 0 153990 800
rect 156510 0 156566 800
rect 159086 0 159142 800
rect 161662 0 161718 800
rect 164882 0 164938 800
rect 167458 0 167514 800
rect 170034 0 170090 800
rect 173254 0 173310 800
rect 175830 0 175886 800
rect 178406 0 178462 800
rect 180982 0 181038 800
rect 184202 0 184258 800
rect 186778 0 186834 800
rect 189354 0 189410 800
rect 191930 0 191986 800
rect 195150 0 195206 800
rect 197726 0 197782 800
rect 200302 0 200358 800
rect 202878 0 202934 800
rect 206098 0 206154 800
rect 208674 0 208730 800
rect 211250 0 211306 800
rect 214470 0 214526 800
rect 217046 0 217102 800
rect 219622 0 219678 800
rect 222198 0 222254 800
rect 225418 0 225474 800
rect 227994 0 228050 800
rect 230570 0 230626 800
rect 233146 0 233202 800
rect 236366 0 236422 800
rect 238942 0 238998 800
rect 241518 0 241574 800
rect 244738 0 244794 800
rect 247314 0 247370 800
rect 249890 0 249946 800
rect 252466 0 252522 800
rect 255686 0 255742 800
rect 258262 0 258318 800
rect 260838 0 260894 800
rect 263414 0 263470 800
rect 266634 0 266690 800
rect 269210 0 269266 800
rect 271786 0 271842 800
rect 275006 0 275062 800
rect 277582 0 277638 800
rect 280158 0 280214 800
rect 282734 0 282790 800
rect 285954 0 286010 800
rect 288530 0 288586 800
rect 291106 0 291162 800
rect 293682 0 293738 800
rect 296902 0 296958 800
rect 299478 0 299534 800
rect 302054 0 302110 800
rect 304630 0 304686 800
rect 307850 0 307906 800
rect 310426 0 310482 800
rect 313002 0 313058 800
rect 316222 0 316278 800
rect 318798 0 318854 800
rect 321374 0 321430 800
rect 323950 0 324006 800
rect 327170 0 327226 800
rect 329746 0 329802 800
rect 332322 0 332378 800
rect 334898 0 334954 800
rect 338118 0 338174 800
rect 340694 0 340750 800
rect 343270 0 343326 800
rect 346490 0 346546 800
rect 349066 0 349122 800
rect 351642 0 351698 800
rect 354218 0 354274 800
rect 357438 0 357494 800
rect 360014 0 360070 800
rect 362590 0 362646 800
rect 365166 0 365222 800
rect 368386 0 368442 800
rect 370962 0 371018 800
rect 373538 0 373594 800
rect 376758 0 376814 800
rect 379334 0 379390 800
<< obsm2 >>
rect 20 479144 1250 479346
rect 1418 479144 4470 479346
rect 4638 479144 7046 479346
rect 7214 479144 9622 479346
rect 9790 479144 12198 479346
rect 12366 479144 15418 479346
rect 15586 479144 17994 479346
rect 18162 479144 20570 479346
rect 20738 479144 23790 479346
rect 23958 479144 26366 479346
rect 26534 479144 28942 479346
rect 29110 479144 31518 479346
rect 31686 479144 34738 479346
rect 34906 479144 37314 479346
rect 37482 479144 39890 479346
rect 40058 479144 42466 479346
rect 42634 479144 45686 479346
rect 45854 479144 48262 479346
rect 48430 479144 50838 479346
rect 51006 479144 53414 479346
rect 53582 479144 56634 479346
rect 56802 479144 59210 479346
rect 59378 479144 61786 479346
rect 61954 479144 65006 479346
rect 65174 479144 67582 479346
rect 67750 479144 70158 479346
rect 70326 479144 72734 479346
rect 72902 479144 75954 479346
rect 76122 479144 78530 479346
rect 78698 479144 81106 479346
rect 81274 479144 83682 479346
rect 83850 479144 86902 479346
rect 87070 479144 89478 479346
rect 89646 479144 92054 479346
rect 92222 479144 95274 479346
rect 95442 479144 97850 479346
rect 98018 479144 100426 479346
rect 100594 479144 103002 479346
rect 103170 479144 106222 479346
rect 106390 479144 108798 479346
rect 108966 479144 111374 479346
rect 111542 479144 113950 479346
rect 114118 479144 117170 479346
rect 117338 479144 119746 479346
rect 119914 479144 122322 479346
rect 122490 479144 125542 479346
rect 125710 479144 128118 479346
rect 128286 479144 130694 479346
rect 130862 479144 133270 479346
rect 133438 479144 136490 479346
rect 136658 479144 139066 479346
rect 139234 479144 141642 479346
rect 141810 479144 144218 479346
rect 144386 479144 147438 479346
rect 147606 479144 150014 479346
rect 150182 479144 152590 479346
rect 152758 479144 155166 479346
rect 155334 479144 158386 479346
rect 158554 479144 160962 479346
rect 161130 479144 163538 479346
rect 163706 479144 166758 479346
rect 166926 479144 169334 479346
rect 169502 479144 171910 479346
rect 172078 479144 174486 479346
rect 174654 479144 177706 479346
rect 177874 479144 180282 479346
rect 180450 479144 182858 479346
rect 183026 479144 185434 479346
rect 185602 479144 188654 479346
rect 188822 479144 191230 479346
rect 191398 479144 193806 479346
rect 193974 479144 197026 479346
rect 197194 479144 199602 479346
rect 199770 479144 202178 479346
rect 202346 479144 204754 479346
rect 204922 479144 207974 479346
rect 208142 479144 210550 479346
rect 210718 479144 213126 479346
rect 213294 479144 215702 479346
rect 215870 479144 218922 479346
rect 219090 479144 221498 479346
rect 221666 479144 224074 479346
rect 224242 479144 227294 479346
rect 227462 479144 229870 479346
rect 230038 479144 232446 479346
rect 232614 479144 235022 479346
rect 235190 479144 238242 479346
rect 238410 479144 240818 479346
rect 240986 479144 243394 479346
rect 243562 479144 245970 479346
rect 246138 479144 249190 479346
rect 249358 479144 251766 479346
rect 251934 479144 254342 479346
rect 254510 479144 256918 479346
rect 257086 479144 260138 479346
rect 260306 479144 262714 479346
rect 262882 479144 265290 479346
rect 265458 479144 268510 479346
rect 268678 479144 271086 479346
rect 271254 479144 273662 479346
rect 273830 479144 276238 479346
rect 276406 479144 279458 479346
rect 279626 479144 282034 479346
rect 282202 479144 284610 479346
rect 284778 479144 287186 479346
rect 287354 479144 290406 479346
rect 290574 479144 292982 479346
rect 293150 479144 295558 479346
rect 295726 479144 298778 479346
rect 298946 479144 301354 479346
rect 301522 479144 303930 479346
rect 304098 479144 306506 479346
rect 306674 479144 309726 479346
rect 309894 479144 312302 479346
rect 312470 479144 314878 479346
rect 315046 479144 317454 479346
rect 317622 479144 320674 479346
rect 320842 479144 323250 479346
rect 323418 479144 325826 479346
rect 325994 479144 329046 479346
rect 329214 479144 331622 479346
rect 331790 479144 334198 479346
rect 334366 479144 336774 479346
rect 336942 479144 339994 479346
rect 340162 479144 342570 479346
rect 342738 479144 345146 479346
rect 345314 479144 347722 479346
rect 347890 479144 350942 479346
rect 351110 479144 353518 479346
rect 353686 479144 356094 479346
rect 356262 479144 358670 479346
rect 358838 479144 361890 479346
rect 362058 479144 364466 479346
rect 364634 479144 367042 479346
rect 367210 479144 370262 479346
rect 370430 479144 372838 479346
rect 373006 479144 375414 479346
rect 375582 479144 377990 479346
rect 378158 479144 379388 479346
rect 20 856 379388 479144
rect 130 800 2538 856
rect 2706 800 5114 856
rect 5282 800 7690 856
rect 7858 800 10910 856
rect 11078 800 13486 856
rect 13654 800 16062 856
rect 16230 800 18638 856
rect 18806 800 21858 856
rect 22026 800 24434 856
rect 24602 800 27010 856
rect 27178 800 29586 856
rect 29754 800 32806 856
rect 32974 800 35382 856
rect 35550 800 37958 856
rect 38126 800 41178 856
rect 41346 800 43754 856
rect 43922 800 46330 856
rect 46498 800 48906 856
rect 49074 800 52126 856
rect 52294 800 54702 856
rect 54870 800 57278 856
rect 57446 800 59854 856
rect 60022 800 63074 856
rect 63242 800 65650 856
rect 65818 800 68226 856
rect 68394 800 71446 856
rect 71614 800 74022 856
rect 74190 800 76598 856
rect 76766 800 79174 856
rect 79342 800 82394 856
rect 82562 800 84970 856
rect 85138 800 87546 856
rect 87714 800 90122 856
rect 90290 800 93342 856
rect 93510 800 95918 856
rect 96086 800 98494 856
rect 98662 800 101070 856
rect 101238 800 104290 856
rect 104458 800 106866 856
rect 107034 800 109442 856
rect 109610 800 112662 856
rect 112830 800 115238 856
rect 115406 800 117814 856
rect 117982 800 120390 856
rect 120558 800 123610 856
rect 123778 800 126186 856
rect 126354 800 128762 856
rect 128930 800 131338 856
rect 131506 800 134558 856
rect 134726 800 137134 856
rect 137302 800 139710 856
rect 139878 800 142930 856
rect 143098 800 145506 856
rect 145674 800 148082 856
rect 148250 800 150658 856
rect 150826 800 153878 856
rect 154046 800 156454 856
rect 156622 800 159030 856
rect 159198 800 161606 856
rect 161774 800 164826 856
rect 164994 800 167402 856
rect 167570 800 169978 856
rect 170146 800 173198 856
rect 173366 800 175774 856
rect 175942 800 178350 856
rect 178518 800 180926 856
rect 181094 800 184146 856
rect 184314 800 186722 856
rect 186890 800 189298 856
rect 189466 800 191874 856
rect 192042 800 195094 856
rect 195262 800 197670 856
rect 197838 800 200246 856
rect 200414 800 202822 856
rect 202990 800 206042 856
rect 206210 800 208618 856
rect 208786 800 211194 856
rect 211362 800 214414 856
rect 214582 800 216990 856
rect 217158 800 219566 856
rect 219734 800 222142 856
rect 222310 800 225362 856
rect 225530 800 227938 856
rect 228106 800 230514 856
rect 230682 800 233090 856
rect 233258 800 236310 856
rect 236478 800 238886 856
rect 239054 800 241462 856
rect 241630 800 244682 856
rect 244850 800 247258 856
rect 247426 800 249834 856
rect 250002 800 252410 856
rect 252578 800 255630 856
rect 255798 800 258206 856
rect 258374 800 260782 856
rect 260950 800 263358 856
rect 263526 800 266578 856
rect 266746 800 269154 856
rect 269322 800 271730 856
rect 271898 800 274950 856
rect 275118 800 277526 856
rect 277694 800 280102 856
rect 280270 800 282678 856
rect 282846 800 285898 856
rect 286066 800 288474 856
rect 288642 800 291050 856
rect 291218 800 293626 856
rect 293794 800 296846 856
rect 297014 800 299422 856
rect 299590 800 301998 856
rect 302166 800 304574 856
rect 304742 800 307794 856
rect 307962 800 310370 856
rect 310538 800 312946 856
rect 313114 800 316166 856
rect 316334 800 318742 856
rect 318910 800 321318 856
rect 321486 800 323894 856
rect 324062 800 327114 856
rect 327282 800 329690 856
rect 329858 800 332266 856
rect 332434 800 334842 856
rect 335010 800 338062 856
rect 338230 800 340638 856
rect 340806 800 343214 856
rect 343382 800 346434 856
rect 346602 800 349010 856
rect 349178 800 351586 856
rect 351754 800 354162 856
rect 354330 800 357382 856
rect 357550 800 359958 856
rect 360126 800 362534 856
rect 362702 800 365110 856
rect 365278 800 368330 856
rect 368498 800 370906 856
rect 371074 800 373482 856
rect 373650 800 376702 856
rect 376870 800 379278 856
<< metal3 >>
rect 0 478728 800 478848
rect 379200 478048 380000 478168
rect 0 476008 800 476128
rect 379200 475328 380000 475448
rect 0 473288 800 473408
rect 379200 472608 380000 472728
rect 0 469888 800 470008
rect 379200 469888 380000 470008
rect 0 467168 800 467288
rect 379200 466488 380000 466608
rect 0 464448 800 464568
rect 379200 463768 380000 463888
rect 0 461048 800 461168
rect 379200 461048 380000 461168
rect 0 458328 800 458448
rect 379200 457648 380000 457768
rect 0 455608 800 455728
rect 379200 454928 380000 455048
rect 0 452888 800 453008
rect 379200 452208 380000 452328
rect 0 449488 800 449608
rect 379200 449488 380000 449608
rect 0 446768 800 446888
rect 379200 446088 380000 446208
rect 0 444048 800 444168
rect 379200 443368 380000 443488
rect 0 441328 800 441448
rect 379200 440648 380000 440768
rect 0 437928 800 438048
rect 379200 437928 380000 438048
rect 0 435208 800 435328
rect 379200 434528 380000 434648
rect 0 432488 800 432608
rect 379200 431808 380000 431928
rect 0 429088 800 429208
rect 379200 429088 380000 429208
rect 0 426368 800 426488
rect 379200 426368 380000 426488
rect 0 423648 800 423768
rect 379200 422968 380000 423088
rect 0 420928 800 421048
rect 379200 420248 380000 420368
rect 0 417528 800 417648
rect 379200 417528 380000 417648
rect 0 414808 800 414928
rect 379200 414128 380000 414248
rect 0 412088 800 412208
rect 379200 411408 380000 411528
rect 0 409368 800 409488
rect 379200 408688 380000 408808
rect 0 405968 800 406088
rect 379200 405968 380000 406088
rect 0 403248 800 403368
rect 379200 402568 380000 402688
rect 0 400528 800 400648
rect 379200 399848 380000 399968
rect 0 397808 800 397928
rect 379200 397128 380000 397248
rect 0 394408 800 394528
rect 379200 394408 380000 394528
rect 0 391688 800 391808
rect 379200 391008 380000 391128
rect 0 388968 800 389088
rect 379200 388288 380000 388408
rect 0 385568 800 385688
rect 379200 385568 380000 385688
rect 0 382848 800 382968
rect 379200 382168 380000 382288
rect 0 380128 800 380248
rect 379200 379448 380000 379568
rect 0 377408 800 377528
rect 379200 376728 380000 376848
rect 0 374008 800 374128
rect 379200 374008 380000 374128
rect 0 371288 800 371408
rect 379200 370608 380000 370728
rect 0 368568 800 368688
rect 379200 367888 380000 368008
rect 0 365848 800 365968
rect 379200 365168 380000 365288
rect 0 362448 800 362568
rect 379200 362448 380000 362568
rect 0 359728 800 359848
rect 379200 359048 380000 359168
rect 0 357008 800 357128
rect 379200 356328 380000 356448
rect 0 353608 800 353728
rect 379200 353608 380000 353728
rect 0 350888 800 351008
rect 379200 350208 380000 350328
rect 0 348168 800 348288
rect 379200 347488 380000 347608
rect 0 345448 800 345568
rect 379200 344768 380000 344888
rect 0 342048 800 342168
rect 379200 342048 380000 342168
rect 0 339328 800 339448
rect 379200 338648 380000 338768
rect 0 336608 800 336728
rect 379200 335928 380000 336048
rect 0 333888 800 334008
rect 379200 333208 380000 333328
rect 0 330488 800 330608
rect 379200 330488 380000 330608
rect 0 327768 800 327888
rect 379200 327088 380000 327208
rect 0 325048 800 325168
rect 379200 324368 380000 324488
rect 0 321648 800 321768
rect 379200 321648 380000 321768
rect 0 318928 800 319048
rect 379200 318928 380000 319048
rect 0 316208 800 316328
rect 379200 315528 380000 315648
rect 0 313488 800 313608
rect 379200 312808 380000 312928
rect 0 310088 800 310208
rect 379200 310088 380000 310208
rect 0 307368 800 307488
rect 379200 306688 380000 306808
rect 0 304648 800 304768
rect 379200 303968 380000 304088
rect 0 301928 800 302048
rect 379200 301248 380000 301368
rect 0 298528 800 298648
rect 379200 298528 380000 298648
rect 0 295808 800 295928
rect 379200 295128 380000 295248
rect 0 293088 800 293208
rect 379200 292408 380000 292528
rect 0 290368 800 290488
rect 379200 289688 380000 289808
rect 0 286968 800 287088
rect 379200 286968 380000 287088
rect 0 284248 800 284368
rect 379200 283568 380000 283688
rect 0 281528 800 281648
rect 379200 280848 380000 280968
rect 0 278128 800 278248
rect 379200 278128 380000 278248
rect 0 275408 800 275528
rect 379200 274728 380000 274848
rect 0 272688 800 272808
rect 379200 272008 380000 272128
rect 0 269968 800 270088
rect 379200 269288 380000 269408
rect 0 266568 800 266688
rect 379200 266568 380000 266688
rect 0 263848 800 263968
rect 379200 263168 380000 263288
rect 0 261128 800 261248
rect 379200 260448 380000 260568
rect 0 258408 800 258528
rect 379200 257728 380000 257848
rect 0 255008 800 255128
rect 379200 255008 380000 255128
rect 0 252288 800 252408
rect 379200 251608 380000 251728
rect 0 249568 800 249688
rect 379200 248888 380000 249008
rect 0 246168 800 246288
rect 379200 246168 380000 246288
rect 0 243448 800 243568
rect 379200 242768 380000 242888
rect 0 240728 800 240848
rect 379200 240048 380000 240168
rect 0 238008 800 238128
rect 379200 237328 380000 237448
rect 0 234608 800 234728
rect 379200 234608 380000 234728
rect 0 231888 800 232008
rect 379200 231208 380000 231328
rect 0 229168 800 229288
rect 379200 228488 380000 228608
rect 0 226448 800 226568
rect 379200 225768 380000 225888
rect 0 223048 800 223168
rect 379200 223048 380000 223168
rect 0 220328 800 220448
rect 379200 219648 380000 219768
rect 0 217608 800 217728
rect 379200 216928 380000 217048
rect 0 214208 800 214328
rect 379200 214208 380000 214328
rect 0 211488 800 211608
rect 379200 211488 380000 211608
rect 0 208768 800 208888
rect 379200 208088 380000 208208
rect 0 206048 800 206168
rect 379200 205368 380000 205488
rect 0 202648 800 202768
rect 379200 202648 380000 202768
rect 0 199928 800 200048
rect 379200 199248 380000 199368
rect 0 197208 800 197328
rect 379200 196528 380000 196648
rect 0 194488 800 194608
rect 379200 193808 380000 193928
rect 0 191088 800 191208
rect 379200 191088 380000 191208
rect 0 188368 800 188488
rect 379200 187688 380000 187808
rect 0 185648 800 185768
rect 379200 184968 380000 185088
rect 0 182928 800 183048
rect 379200 182248 380000 182368
rect 0 179528 800 179648
rect 379200 179528 380000 179648
rect 0 176808 800 176928
rect 379200 176128 380000 176248
rect 0 174088 800 174208
rect 379200 173408 380000 173528
rect 0 170688 800 170808
rect 379200 170688 380000 170808
rect 0 167968 800 168088
rect 379200 167288 380000 167408
rect 0 165248 800 165368
rect 379200 164568 380000 164688
rect 0 162528 800 162648
rect 379200 161848 380000 161968
rect 0 159128 800 159248
rect 379200 159128 380000 159248
rect 0 156408 800 156528
rect 379200 155728 380000 155848
rect 0 153688 800 153808
rect 379200 153008 380000 153128
rect 0 150968 800 151088
rect 379200 150288 380000 150408
rect 0 147568 800 147688
rect 379200 147568 380000 147688
rect 0 144848 800 144968
rect 379200 144168 380000 144288
rect 0 142128 800 142248
rect 379200 141448 380000 141568
rect 0 138728 800 138848
rect 379200 138728 380000 138848
rect 0 136008 800 136128
rect 379200 135328 380000 135448
rect 0 133288 800 133408
rect 379200 132608 380000 132728
rect 0 130568 800 130688
rect 379200 129888 380000 130008
rect 0 127168 800 127288
rect 379200 127168 380000 127288
rect 0 124448 800 124568
rect 379200 123768 380000 123888
rect 0 121728 800 121848
rect 379200 121048 380000 121168
rect 0 119008 800 119128
rect 379200 118328 380000 118448
rect 0 115608 800 115728
rect 379200 115608 380000 115728
rect 0 112888 800 113008
rect 379200 112208 380000 112328
rect 0 110168 800 110288
rect 379200 109488 380000 109608
rect 0 106768 800 106888
rect 379200 106768 380000 106888
rect 0 104048 800 104168
rect 379200 104048 380000 104168
rect 0 101328 800 101448
rect 379200 100648 380000 100768
rect 0 98608 800 98728
rect 379200 97928 380000 98048
rect 0 95208 800 95328
rect 379200 95208 380000 95328
rect 0 92488 800 92608
rect 379200 91808 380000 91928
rect 0 89768 800 89888
rect 379200 89088 380000 89208
rect 0 87048 800 87168
rect 379200 86368 380000 86488
rect 0 83648 800 83768
rect 379200 83648 380000 83768
rect 0 80928 800 81048
rect 379200 80248 380000 80368
rect 0 78208 800 78328
rect 379200 77528 380000 77648
rect 0 75488 800 75608
rect 379200 74808 380000 74928
rect 0 72088 800 72208
rect 379200 72088 380000 72208
rect 0 69368 800 69488
rect 379200 68688 380000 68808
rect 0 66648 800 66768
rect 379200 65968 380000 66088
rect 0 63248 800 63368
rect 379200 63248 380000 63368
rect 0 60528 800 60648
rect 379200 59848 380000 59968
rect 0 57808 800 57928
rect 379200 57128 380000 57248
rect 0 55088 800 55208
rect 379200 54408 380000 54528
rect 0 51688 800 51808
rect 379200 51688 380000 51808
rect 0 48968 800 49088
rect 379200 48288 380000 48408
rect 0 46248 800 46368
rect 379200 45568 380000 45688
rect 0 43528 800 43648
rect 379200 42848 380000 42968
rect 0 40128 800 40248
rect 379200 40128 380000 40248
rect 0 37408 800 37528
rect 379200 36728 380000 36848
rect 0 34688 800 34808
rect 379200 34008 380000 34128
rect 0 31288 800 31408
rect 379200 31288 380000 31408
rect 0 28568 800 28688
rect 379200 27888 380000 28008
rect 0 25848 800 25968
rect 379200 25168 380000 25288
rect 0 23128 800 23248
rect 379200 22448 380000 22568
rect 0 19728 800 19848
rect 379200 19728 380000 19848
rect 0 17008 800 17128
rect 379200 16328 380000 16448
rect 0 14288 800 14408
rect 379200 13608 380000 13728
rect 0 11568 800 11688
rect 379200 10888 380000 11008
rect 0 8168 800 8288
rect 379200 8168 380000 8288
rect 0 5448 800 5568
rect 379200 4768 380000 4888
rect 0 2728 800 2848
rect 379200 2048 380000 2168
<< obsm3 >>
rect 880 478648 379200 478821
rect 800 478248 379200 478648
rect 800 477968 379120 478248
rect 800 476208 379200 477968
rect 880 475928 379200 476208
rect 800 475528 379200 475928
rect 800 475248 379120 475528
rect 800 473488 379200 475248
rect 880 473208 379200 473488
rect 800 472808 379200 473208
rect 800 472528 379120 472808
rect 800 470088 379200 472528
rect 880 469808 379120 470088
rect 800 467368 379200 469808
rect 880 467088 379200 467368
rect 800 466688 379200 467088
rect 800 466408 379120 466688
rect 800 464648 379200 466408
rect 880 464368 379200 464648
rect 800 463968 379200 464368
rect 800 463688 379120 463968
rect 800 461248 379200 463688
rect 880 460968 379120 461248
rect 800 458528 379200 460968
rect 880 458248 379200 458528
rect 800 457848 379200 458248
rect 800 457568 379120 457848
rect 800 455808 379200 457568
rect 880 455528 379200 455808
rect 800 455128 379200 455528
rect 800 454848 379120 455128
rect 800 453088 379200 454848
rect 880 452808 379200 453088
rect 800 452408 379200 452808
rect 800 452128 379120 452408
rect 800 449688 379200 452128
rect 880 449408 379120 449688
rect 800 446968 379200 449408
rect 880 446688 379200 446968
rect 800 446288 379200 446688
rect 800 446008 379120 446288
rect 800 444248 379200 446008
rect 880 443968 379200 444248
rect 800 443568 379200 443968
rect 800 443288 379120 443568
rect 800 441528 379200 443288
rect 880 441248 379200 441528
rect 800 440848 379200 441248
rect 800 440568 379120 440848
rect 800 438128 379200 440568
rect 880 437848 379120 438128
rect 800 435408 379200 437848
rect 880 435128 379200 435408
rect 800 434728 379200 435128
rect 800 434448 379120 434728
rect 800 432688 379200 434448
rect 880 432408 379200 432688
rect 800 432008 379200 432408
rect 800 431728 379120 432008
rect 800 429288 379200 431728
rect 880 429008 379120 429288
rect 800 426568 379200 429008
rect 880 426288 379120 426568
rect 800 423848 379200 426288
rect 880 423568 379200 423848
rect 800 423168 379200 423568
rect 800 422888 379120 423168
rect 800 421128 379200 422888
rect 880 420848 379200 421128
rect 800 420448 379200 420848
rect 800 420168 379120 420448
rect 800 417728 379200 420168
rect 880 417448 379120 417728
rect 800 415008 379200 417448
rect 880 414728 379200 415008
rect 800 414328 379200 414728
rect 800 414048 379120 414328
rect 800 412288 379200 414048
rect 880 412008 379200 412288
rect 800 411608 379200 412008
rect 800 411328 379120 411608
rect 800 409568 379200 411328
rect 880 409288 379200 409568
rect 800 408888 379200 409288
rect 800 408608 379120 408888
rect 800 406168 379200 408608
rect 880 405888 379120 406168
rect 800 403448 379200 405888
rect 880 403168 379200 403448
rect 800 402768 379200 403168
rect 800 402488 379120 402768
rect 800 400728 379200 402488
rect 880 400448 379200 400728
rect 800 400048 379200 400448
rect 800 399768 379120 400048
rect 800 398008 379200 399768
rect 880 397728 379200 398008
rect 800 397328 379200 397728
rect 800 397048 379120 397328
rect 800 394608 379200 397048
rect 880 394328 379120 394608
rect 800 391888 379200 394328
rect 880 391608 379200 391888
rect 800 391208 379200 391608
rect 800 390928 379120 391208
rect 800 389168 379200 390928
rect 880 388888 379200 389168
rect 800 388488 379200 388888
rect 800 388208 379120 388488
rect 800 385768 379200 388208
rect 880 385488 379120 385768
rect 800 383048 379200 385488
rect 880 382768 379200 383048
rect 800 382368 379200 382768
rect 800 382088 379120 382368
rect 800 380328 379200 382088
rect 880 380048 379200 380328
rect 800 379648 379200 380048
rect 800 379368 379120 379648
rect 800 377608 379200 379368
rect 880 377328 379200 377608
rect 800 376928 379200 377328
rect 800 376648 379120 376928
rect 800 374208 379200 376648
rect 880 373928 379120 374208
rect 800 371488 379200 373928
rect 880 371208 379200 371488
rect 800 370808 379200 371208
rect 800 370528 379120 370808
rect 800 368768 379200 370528
rect 880 368488 379200 368768
rect 800 368088 379200 368488
rect 800 367808 379120 368088
rect 800 366048 379200 367808
rect 880 365768 379200 366048
rect 800 365368 379200 365768
rect 800 365088 379120 365368
rect 800 362648 379200 365088
rect 880 362368 379120 362648
rect 800 359928 379200 362368
rect 880 359648 379200 359928
rect 800 359248 379200 359648
rect 800 358968 379120 359248
rect 800 357208 379200 358968
rect 880 356928 379200 357208
rect 800 356528 379200 356928
rect 800 356248 379120 356528
rect 800 353808 379200 356248
rect 880 353528 379120 353808
rect 800 351088 379200 353528
rect 880 350808 379200 351088
rect 800 350408 379200 350808
rect 800 350128 379120 350408
rect 800 348368 379200 350128
rect 880 348088 379200 348368
rect 800 347688 379200 348088
rect 800 347408 379120 347688
rect 800 345648 379200 347408
rect 880 345368 379200 345648
rect 800 344968 379200 345368
rect 800 344688 379120 344968
rect 800 342248 379200 344688
rect 880 341968 379120 342248
rect 800 339528 379200 341968
rect 880 339248 379200 339528
rect 800 338848 379200 339248
rect 800 338568 379120 338848
rect 800 336808 379200 338568
rect 880 336528 379200 336808
rect 800 336128 379200 336528
rect 800 335848 379120 336128
rect 800 334088 379200 335848
rect 880 333808 379200 334088
rect 800 333408 379200 333808
rect 800 333128 379120 333408
rect 800 330688 379200 333128
rect 880 330408 379120 330688
rect 800 327968 379200 330408
rect 880 327688 379200 327968
rect 800 327288 379200 327688
rect 800 327008 379120 327288
rect 800 325248 379200 327008
rect 880 324968 379200 325248
rect 800 324568 379200 324968
rect 800 324288 379120 324568
rect 800 321848 379200 324288
rect 880 321568 379120 321848
rect 800 319128 379200 321568
rect 880 318848 379120 319128
rect 800 316408 379200 318848
rect 880 316128 379200 316408
rect 800 315728 379200 316128
rect 800 315448 379120 315728
rect 800 313688 379200 315448
rect 880 313408 379200 313688
rect 800 313008 379200 313408
rect 800 312728 379120 313008
rect 800 310288 379200 312728
rect 880 310008 379120 310288
rect 800 307568 379200 310008
rect 880 307288 379200 307568
rect 800 306888 379200 307288
rect 800 306608 379120 306888
rect 800 304848 379200 306608
rect 880 304568 379200 304848
rect 800 304168 379200 304568
rect 800 303888 379120 304168
rect 800 302128 379200 303888
rect 880 301848 379200 302128
rect 800 301448 379200 301848
rect 800 301168 379120 301448
rect 800 298728 379200 301168
rect 880 298448 379120 298728
rect 800 296008 379200 298448
rect 880 295728 379200 296008
rect 800 295328 379200 295728
rect 800 295048 379120 295328
rect 800 293288 379200 295048
rect 880 293008 379200 293288
rect 800 292608 379200 293008
rect 800 292328 379120 292608
rect 800 290568 379200 292328
rect 880 290288 379200 290568
rect 800 289888 379200 290288
rect 800 289608 379120 289888
rect 800 287168 379200 289608
rect 880 286888 379120 287168
rect 800 284448 379200 286888
rect 880 284168 379200 284448
rect 800 283768 379200 284168
rect 800 283488 379120 283768
rect 800 281728 379200 283488
rect 880 281448 379200 281728
rect 800 281048 379200 281448
rect 800 280768 379120 281048
rect 800 278328 379200 280768
rect 880 278048 379120 278328
rect 800 275608 379200 278048
rect 880 275328 379200 275608
rect 800 274928 379200 275328
rect 800 274648 379120 274928
rect 800 272888 379200 274648
rect 880 272608 379200 272888
rect 800 272208 379200 272608
rect 800 271928 379120 272208
rect 800 270168 379200 271928
rect 880 269888 379200 270168
rect 800 269488 379200 269888
rect 800 269208 379120 269488
rect 800 266768 379200 269208
rect 880 266488 379120 266768
rect 800 264048 379200 266488
rect 880 263768 379200 264048
rect 800 263368 379200 263768
rect 800 263088 379120 263368
rect 800 261328 379200 263088
rect 880 261048 379200 261328
rect 800 260648 379200 261048
rect 800 260368 379120 260648
rect 800 258608 379200 260368
rect 880 258328 379200 258608
rect 800 257928 379200 258328
rect 800 257648 379120 257928
rect 800 255208 379200 257648
rect 880 254928 379120 255208
rect 800 252488 379200 254928
rect 880 252208 379200 252488
rect 800 251808 379200 252208
rect 800 251528 379120 251808
rect 800 249768 379200 251528
rect 880 249488 379200 249768
rect 800 249088 379200 249488
rect 800 248808 379120 249088
rect 800 246368 379200 248808
rect 880 246088 379120 246368
rect 800 243648 379200 246088
rect 880 243368 379200 243648
rect 800 242968 379200 243368
rect 800 242688 379120 242968
rect 800 240928 379200 242688
rect 880 240648 379200 240928
rect 800 240248 379200 240648
rect 800 239968 379120 240248
rect 800 238208 379200 239968
rect 880 237928 379200 238208
rect 800 237528 379200 237928
rect 800 237248 379120 237528
rect 800 234808 379200 237248
rect 880 234528 379120 234808
rect 800 232088 379200 234528
rect 880 231808 379200 232088
rect 800 231408 379200 231808
rect 800 231128 379120 231408
rect 800 229368 379200 231128
rect 880 229088 379200 229368
rect 800 228688 379200 229088
rect 800 228408 379120 228688
rect 800 226648 379200 228408
rect 880 226368 379200 226648
rect 800 225968 379200 226368
rect 800 225688 379120 225968
rect 800 223248 379200 225688
rect 880 222968 379120 223248
rect 800 220528 379200 222968
rect 880 220248 379200 220528
rect 800 219848 379200 220248
rect 800 219568 379120 219848
rect 800 217808 379200 219568
rect 880 217528 379200 217808
rect 800 217128 379200 217528
rect 800 216848 379120 217128
rect 800 214408 379200 216848
rect 880 214128 379120 214408
rect 800 211688 379200 214128
rect 880 211408 379120 211688
rect 800 208968 379200 211408
rect 880 208688 379200 208968
rect 800 208288 379200 208688
rect 800 208008 379120 208288
rect 800 206248 379200 208008
rect 880 205968 379200 206248
rect 800 205568 379200 205968
rect 800 205288 379120 205568
rect 800 202848 379200 205288
rect 880 202568 379120 202848
rect 800 200128 379200 202568
rect 880 199848 379200 200128
rect 800 199448 379200 199848
rect 800 199168 379120 199448
rect 800 197408 379200 199168
rect 880 197128 379200 197408
rect 800 196728 379200 197128
rect 800 196448 379120 196728
rect 800 194688 379200 196448
rect 880 194408 379200 194688
rect 800 194008 379200 194408
rect 800 193728 379120 194008
rect 800 191288 379200 193728
rect 880 191008 379120 191288
rect 800 188568 379200 191008
rect 880 188288 379200 188568
rect 800 187888 379200 188288
rect 800 187608 379120 187888
rect 800 185848 379200 187608
rect 880 185568 379200 185848
rect 800 185168 379200 185568
rect 800 184888 379120 185168
rect 800 183128 379200 184888
rect 880 182848 379200 183128
rect 800 182448 379200 182848
rect 800 182168 379120 182448
rect 800 179728 379200 182168
rect 880 179448 379120 179728
rect 800 177008 379200 179448
rect 880 176728 379200 177008
rect 800 176328 379200 176728
rect 800 176048 379120 176328
rect 800 174288 379200 176048
rect 880 174008 379200 174288
rect 800 173608 379200 174008
rect 800 173328 379120 173608
rect 800 170888 379200 173328
rect 880 170608 379120 170888
rect 800 168168 379200 170608
rect 880 167888 379200 168168
rect 800 167488 379200 167888
rect 800 167208 379120 167488
rect 800 165448 379200 167208
rect 880 165168 379200 165448
rect 800 164768 379200 165168
rect 800 164488 379120 164768
rect 800 162728 379200 164488
rect 880 162448 379200 162728
rect 800 162048 379200 162448
rect 800 161768 379120 162048
rect 800 159328 379200 161768
rect 880 159048 379120 159328
rect 800 156608 379200 159048
rect 880 156328 379200 156608
rect 800 155928 379200 156328
rect 800 155648 379120 155928
rect 800 153888 379200 155648
rect 880 153608 379200 153888
rect 800 153208 379200 153608
rect 800 152928 379120 153208
rect 800 151168 379200 152928
rect 880 150888 379200 151168
rect 800 150488 379200 150888
rect 800 150208 379120 150488
rect 800 147768 379200 150208
rect 880 147488 379120 147768
rect 800 145048 379200 147488
rect 880 144768 379200 145048
rect 800 144368 379200 144768
rect 800 144088 379120 144368
rect 800 142328 379200 144088
rect 880 142048 379200 142328
rect 800 141648 379200 142048
rect 800 141368 379120 141648
rect 800 138928 379200 141368
rect 880 138648 379120 138928
rect 800 136208 379200 138648
rect 880 135928 379200 136208
rect 800 135528 379200 135928
rect 800 135248 379120 135528
rect 800 133488 379200 135248
rect 880 133208 379200 133488
rect 800 132808 379200 133208
rect 800 132528 379120 132808
rect 800 130768 379200 132528
rect 880 130488 379200 130768
rect 800 130088 379200 130488
rect 800 129808 379120 130088
rect 800 127368 379200 129808
rect 880 127088 379120 127368
rect 800 124648 379200 127088
rect 880 124368 379200 124648
rect 800 123968 379200 124368
rect 800 123688 379120 123968
rect 800 121928 379200 123688
rect 880 121648 379200 121928
rect 800 121248 379200 121648
rect 800 120968 379120 121248
rect 800 119208 379200 120968
rect 880 118928 379200 119208
rect 800 118528 379200 118928
rect 800 118248 379120 118528
rect 800 115808 379200 118248
rect 880 115528 379120 115808
rect 800 113088 379200 115528
rect 880 112808 379200 113088
rect 800 112408 379200 112808
rect 800 112128 379120 112408
rect 800 110368 379200 112128
rect 880 110088 379200 110368
rect 800 109688 379200 110088
rect 800 109408 379120 109688
rect 800 106968 379200 109408
rect 880 106688 379120 106968
rect 800 104248 379200 106688
rect 880 103968 379120 104248
rect 800 101528 379200 103968
rect 880 101248 379200 101528
rect 800 100848 379200 101248
rect 800 100568 379120 100848
rect 800 98808 379200 100568
rect 880 98528 379200 98808
rect 800 98128 379200 98528
rect 800 97848 379120 98128
rect 800 95408 379200 97848
rect 880 95128 379120 95408
rect 800 92688 379200 95128
rect 880 92408 379200 92688
rect 800 92008 379200 92408
rect 800 91728 379120 92008
rect 800 89968 379200 91728
rect 880 89688 379200 89968
rect 800 89288 379200 89688
rect 800 89008 379120 89288
rect 800 87248 379200 89008
rect 880 86968 379200 87248
rect 800 86568 379200 86968
rect 800 86288 379120 86568
rect 800 83848 379200 86288
rect 880 83568 379120 83848
rect 800 81128 379200 83568
rect 880 80848 379200 81128
rect 800 80448 379200 80848
rect 800 80168 379120 80448
rect 800 78408 379200 80168
rect 880 78128 379200 78408
rect 800 77728 379200 78128
rect 800 77448 379120 77728
rect 800 75688 379200 77448
rect 880 75408 379200 75688
rect 800 75008 379200 75408
rect 800 74728 379120 75008
rect 800 72288 379200 74728
rect 880 72008 379120 72288
rect 800 69568 379200 72008
rect 880 69288 379200 69568
rect 800 68888 379200 69288
rect 800 68608 379120 68888
rect 800 66848 379200 68608
rect 880 66568 379200 66848
rect 800 66168 379200 66568
rect 800 65888 379120 66168
rect 800 63448 379200 65888
rect 880 63168 379120 63448
rect 800 60728 379200 63168
rect 880 60448 379200 60728
rect 800 60048 379200 60448
rect 800 59768 379120 60048
rect 800 58008 379200 59768
rect 880 57728 379200 58008
rect 800 57328 379200 57728
rect 800 57048 379120 57328
rect 800 55288 379200 57048
rect 880 55008 379200 55288
rect 800 54608 379200 55008
rect 800 54328 379120 54608
rect 800 51888 379200 54328
rect 880 51608 379120 51888
rect 800 49168 379200 51608
rect 880 48888 379200 49168
rect 800 48488 379200 48888
rect 800 48208 379120 48488
rect 800 46448 379200 48208
rect 880 46168 379200 46448
rect 800 45768 379200 46168
rect 800 45488 379120 45768
rect 800 43728 379200 45488
rect 880 43448 379200 43728
rect 800 43048 379200 43448
rect 800 42768 379120 43048
rect 800 40328 379200 42768
rect 880 40048 379120 40328
rect 800 37608 379200 40048
rect 880 37328 379200 37608
rect 800 36928 379200 37328
rect 800 36648 379120 36928
rect 800 34888 379200 36648
rect 880 34608 379200 34888
rect 800 34208 379200 34608
rect 800 33928 379120 34208
rect 800 31488 379200 33928
rect 880 31208 379120 31488
rect 800 28768 379200 31208
rect 880 28488 379200 28768
rect 800 28088 379200 28488
rect 800 27808 379120 28088
rect 800 26048 379200 27808
rect 880 25768 379200 26048
rect 800 25368 379200 25768
rect 800 25088 379120 25368
rect 800 23328 379200 25088
rect 880 23048 379200 23328
rect 800 22648 379200 23048
rect 800 22368 379120 22648
rect 800 19928 379200 22368
rect 880 19648 379120 19928
rect 800 17208 379200 19648
rect 880 16928 379200 17208
rect 800 16528 379200 16928
rect 800 16248 379120 16528
rect 800 14488 379200 16248
rect 880 14208 379200 14488
rect 800 13808 379200 14208
rect 800 13528 379120 13808
rect 800 11768 379200 13528
rect 880 11488 379200 11768
rect 800 11088 379200 11488
rect 800 10808 379120 11088
rect 800 8368 379200 10808
rect 880 8088 379120 8368
rect 800 5648 379200 8088
rect 880 5368 379200 5648
rect 800 4968 379200 5368
rect 800 4688 379120 4968
rect 800 2928 379200 4688
rect 880 2648 379200 2928
rect 800 2248 379200 2648
rect 800 2075 379120 2248
<< metal4 >>
rect 4208 2128 4528 477680
rect 19568 2128 19888 477680
rect 34928 2128 35248 477680
rect 50288 2128 50608 477680
rect 65648 2128 65968 477680
rect 81008 2128 81328 477680
rect 96368 2128 96688 477680
rect 111728 2128 112048 477680
rect 127088 2128 127408 477680
rect 142448 2128 142768 477680
rect 157808 2128 158128 477680
rect 173168 2128 173488 477680
rect 188528 2128 188848 477680
rect 203888 2128 204208 477680
rect 219248 2128 219568 477680
rect 234608 2128 234928 477680
rect 249968 2128 250288 477680
rect 265328 2128 265648 477680
rect 280688 2128 281008 477680
rect 296048 2128 296368 477680
rect 311408 2128 311728 477680
rect 326768 2128 327088 477680
rect 342128 2128 342448 477680
rect 357488 2128 357808 477680
rect 372848 2128 373168 477680
<< obsm4 >>
rect 234475 196555 234528 198933
rect 235008 196555 235093 198933
<< labels >>
rlabel metal3 s 379200 31288 380000 31408 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 379200 237328 380000 237448 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 97906 479200 97962 480000 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 379200 330488 380000 330608 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 76010 479200 76066 480000 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 379200 461048 380000 461168 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 111430 479200 111486 480000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 61842 479200 61898 480000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 83738 479200 83794 480000 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 379200 367888 380000 368008 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 449488 800 449608 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 221554 479200 221610 480000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 70214 479200 70270 480000 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 147494 479200 147550 480000 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 0 359728 800 359848 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 243450 479200 243506 480000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 202234 479200 202290 480000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 379200 333208 380000 333328 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 379200 8168 380000 8288 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 356150 479200 356206 480000 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 379200 97928 380000 98048 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 379200 301248 380000 301368 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 243448 800 243568 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 158442 479200 158498 480000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 284248 800 284368 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 379200 199248 380000 199368 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 379200 191088 380000 191208 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 208030 479200 208086 480000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 103058 479200 103114 480000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 310426 0 310482 800 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 28998 479200 29054 480000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 379200 202648 380000 202768 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 io_oeb[16]
port 46 nsew signal output
rlabel metal3 s 0 435208 800 435328 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 0 444048 800 444168 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 282734 0 282790 800 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 31574 479200 31630 480000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 246026 479200 246082 480000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 379200 223048 380000 223168 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 379200 475328 380000 475448 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 342048 800 342168 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 4526 479200 4582 480000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 213182 479200 213238 480000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 379200 365168 380000 365288 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 379200 420248 380000 420368 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 260838 0 260894 800 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 385568 800 385688 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 9678 479200 9734 480000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 452888 800 453008 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 34794 479200 34850 480000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 238008 800 238128 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 186778 0 186834 800 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 321648 800 321768 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 279514 479200 279570 480000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 211250 0 211306 800 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 260194 479200 260250 480000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 364522 479200 364578 480000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 0 310088 800 310208 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 0 478728 800 478848 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 0 429088 800 429208 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 353574 479200 353630 480000 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 0 199928 800 200048 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 379200 449488 380000 449608 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 0 142128 800 142248 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 379200 382168 380000 382288 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 379200 144168 380000 144288 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 379200 327088 380000 327208 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 379200 434528 380000 434648 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 379200 385568 380000 385688 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 321374 0 321430 800 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 423648 800 423768 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 379200 19728 380000 19848 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 233146 0 233202 800 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 379200 91808 380000 91928 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 298528 800 298648 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 39946 479200 40002 480000 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 379200 42848 380000 42968 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 379200 286968 380000 287088 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 361946 479200 362002 480000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 379200 429088 380000 429208 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 379334 0 379390 800 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 379200 374008 380000 374128 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 375470 479200 375526 480000 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 379200 338648 380000 338768 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 37370 479200 37426 480000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 376758 0 376814 800 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 0 214208 800 214328 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 379200 86368 380000 86488 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 379200 315528 380000 315648 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 169390 479200 169446 480000 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 128174 479200 128230 480000 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 0 426368 800 426488 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 379200 219648 380000 219768 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 290462 479200 290518 480000 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 379200 266568 380000 266688 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 379200 167288 380000 167408 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 141698 479200 141754 480000 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 23846 479200 23902 480000 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 379200 443368 380000 443488 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 330488 800 330608 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 379200 318928 380000 319048 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 379200 89088 380000 89208 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 185490 479200 185546 480000 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 379200 159128 380000 159248 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 256974 479200 257030 480000 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 339328 800 339448 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 379200 321648 380000 321768 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 345448 800 345568 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 379200 112208 380000 112328 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 268566 479200 268622 480000 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 125598 479200 125654 480000 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 295614 479200 295670 480000 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 379200 306688 380000 306808 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 316208 800 316328 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 240874 479200 240930 480000 6 la_data_in[120]
port 141 nsew signal input
rlabel metal3 s 379200 27888 380000 28008 6 la_data_in[121]
port 142 nsew signal input
rlabel metal3 s 0 455608 800 455728 6 la_data_in[122]
port 143 nsew signal input
rlabel metal3 s 379200 48288 380000 48408 6 la_data_in[123]
port 144 nsew signal input
rlabel metal3 s 0 473288 800 473408 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 318798 0 318854 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 234608 800 234728 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 370962 0 371018 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 379200 359048 380000 359168 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 379200 228488 380000 228608 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 379200 411408 380000 411528 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 276294 479200 276350 480000 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal3 s 0 441328 800 441448 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 379200 274728 380000 274848 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 379200 129888 380000 130008 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 290368 800 290488 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 379200 394408 380000 394528 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 379200 303968 380000 304088 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 299478 0 299534 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 332322 0 332378 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal3 s 379200 13608 380000 13728 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 108854 479200 108910 480000 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 150070 479200 150126 480000 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 0 365848 800 365968 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 287242 479200 287298 480000 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 367098 479200 367154 480000 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 379200 234608 380000 234728 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 226448 800 226568 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 379200 242768 380000 242888 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 379200 379448 380000 379568 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 95330 479200 95386 480000 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 240728 800 240848 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 280158 0 280214 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 254398 479200 254454 480000 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 la_data_in[50]
port 191 nsew signal input
rlabel metal3 s 0 437928 800 438048 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 358726 479200 358782 480000 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 379200 127168 380000 127288 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 313002 0 313058 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 306562 479200 306618 480000 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 365166 0 365222 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 185648 800 185768 6 la_data_in[5]
port 201 nsew signal input
rlabel metal3 s 0 467168 800 467288 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 379200 150288 380000 150408 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 246168 800 246288 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 379200 454928 380000 455048 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 362590 0 362646 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 0 412088 800 412208 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 130750 479200 130806 480000 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 379200 362448 380000 362568 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 379200 216928 380000 217048 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 379200 153008 380000 153128 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 379200 123768 380000 123888 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 59266 479200 59322 480000 6 la_data_in[72]
port 215 nsew signal input
rlabel metal3 s 379200 36728 380000 36848 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 202878 0 202934 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 379200 324368 380000 324488 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 379200 391008 380000 391128 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 379200 164568 380000 164688 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 379200 179528 380000 179648 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 343270 0 343326 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 379200 182248 380000 182368 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 194488 800 194608 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 309782 479200 309838 480000 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 122378 479200 122434 480000 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 379200 353608 380000 353728 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 220328 800 220448 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 266568 800 266688 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 100482 479200 100538 480000 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 53470 479200 53526 480000 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 199658 479200 199714 480000 6 la_data_in[90]
port 235 nsew signal input
rlabel metal3 s 0 446768 800 446888 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 379200 51688 380000 51808 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 379200 80248 380000 80368 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 0 382848 800 382968 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 379200 248888 380000 249008 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 295808 800 295928 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 275408 800 275528 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 347778 479200 347834 480000 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 0 380128 800 380248 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 379200 205368 380000 205488 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 379200 280848 380000 280968 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 50894 479200 50950 480000 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 275006 0 275062 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 0 348168 800 348288 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 174542 479200 174598 480000 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 210606 479200 210662 480000 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 265346 479200 265402 480000 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 340050 479200 340106 480000 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 133326 479200 133382 480000 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 379200 426368 380000 426488 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 379200 141448 380000 141568 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 159128 800 159248 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 379200 57128 380000 57248 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 26422 479200 26478 480000 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 345202 479200 345258 480000 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 0 350888 800 351008 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 144848 800 144968 6 la_data_out[124]
port 273 nsew signal output
rlabel metal3 s 379200 2048 380000 2168 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 263848 800 263968 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 379200 431808 380000 431928 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 379200 240048 380000 240168 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 379200 260448 380000 260568 6 la_data_out[15]
port 280 nsew signal output
rlabel metal3 s 379200 34008 380000 34128 6 la_data_out[16]
port 281 nsew signal output
rlabel metal3 s 0 469888 800 470008 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 379200 118328 380000 118448 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 281528 800 281648 6 la_data_out[19]
port 284 nsew signal output
rlabel metal3 s 0 464448 800 464568 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 379200 466488 380000 466608 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 232502 479200 232558 480000 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 379200 208088 380000 208208 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 191286 479200 191342 480000 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 379200 246168 380000 246288 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 0 405968 800 406088 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 379200 106768 380000 106888 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 45742 479200 45798 480000 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 197082 479200 197138 480000 6 la_data_out[33]
port 300 nsew signal output
rlabel metal3 s 379200 25168 380000 25288 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 329102 479200 329158 480000 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 327768 800 327888 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 208768 800 208888 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 293038 479200 293094 480000 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 379200 161848 380000 161968 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 117226 479200 117282 480000 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 278128 800 278248 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 236366 0 236422 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 86958 479200 87014 480000 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 72790 479200 72846 480000 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 351642 0 351698 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 379200 54408 380000 54528 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 372894 479200 372950 480000 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 106278 479200 106334 480000 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 206048 800 206168 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 249568 800 249688 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 333888 800 334008 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 379200 263168 380000 263288 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 269968 800 270088 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 379200 251608 380000 251728 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 350998 479200 351054 480000 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 282090 479200 282146 480000 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 161018 479200 161074 480000 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 329746 0 329802 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 0 374008 800 374128 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 379200 278128 380000 278248 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 379200 138728 380000 138848 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 379200 100648 380000 100768 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 200302 0 200358 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 296902 0 296958 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 336830 479200 336886 480000 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 227994 0 228050 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 119802 479200 119858 480000 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 0 414808 800 414928 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 166814 479200 166870 480000 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 208674 0 208730 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 379200 83648 380000 83768 6 la_data_out[75]
port 346 nsew signal output
rlabel metal3 s 379200 16328 380000 16448 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 379200 135328 380000 135448 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 379200 115608 380000 115728 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 0 403248 800 403368 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 48318 479200 48374 480000 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 340694 0 340750 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 18050 479200 18106 480000 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 la_data_out[84]
port 356 nsew signal output
rlabel metal3 s 379200 40128 380000 40248 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 379200 269288 380000 269408 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 188710 479200 188766 480000 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 266634 0 266690 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 177762 479200 177818 480000 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 180338 479200 180394 480000 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 316222 0 316278 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 354218 0 354274 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 314934 479200 314990 480000 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 92110 479200 92166 480000 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 136546 479200 136602 480000 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 327170 0 327226 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal3 s 0 476008 800 476128 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 303986 479200 304042 480000 6 la_data_out[98]
port 371 nsew signal output
rlabel metal3 s 379200 45568 380000 45688 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 222198 0 222254 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 379200 472608 380000 472728 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 0 368568 800 368688 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 312358 479200 312414 480000 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 379200 295128 380000 295248 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 152646 479200 152702 480000 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 370318 479200 370374 480000 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 379200 289688 380000 289808 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 235078 479200 235134 480000 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 284666 479200 284722 480000 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 379200 376728 380000 376848 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 229168 800 229288 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 204810 479200 204866 480000 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 379200 457648 380000 457768 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 379200 214208 380000 214328 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 379200 292408 380000 292528 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 318928 800 319048 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 379200 405968 380000 406088 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 255008 800 255128 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 301928 800 302048 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 346490 0 346546 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 379200 155728 380000 155848 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 379200 344768 380000 344888 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 379200 121048 380000 121168 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 379200 109488 380000 109608 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 379200 452208 380000 452328 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 379200 225768 380000 225888 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 293682 0 293738 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 325882 479200 325938 480000 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 271786 0 271842 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 379200 283568 380000 283688 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 378046 479200 378102 480000 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 331678 479200 331734 480000 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 202648 800 202768 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 78586 479200 78642 480000 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 7102 479200 7158 480000 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 379200 184968 380000 185088 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 379200 298528 380000 298648 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 323950 0 324006 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 379200 399848 380000 399968 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 293088 800 293208 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 342626 479200 342682 480000 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 0 377408 800 377528 6 la_oenb[40]
port 436 nsew signal input
rlabel metal3 s 379200 10888 380000 11008 6 la_oenb[41]
port 437 nsew signal input
rlabel metal3 s 0 458328 800 458448 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 0 371288 800 371408 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 379200 72088 380000 72208 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal3 s 379200 22448 380000 22568 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 379200 176128 380000 176248 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 379200 402568 380000 402688 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 304648 800 304768 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 155222 479200 155278 480000 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 89534 479200 89590 480000 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 217608 800 217728 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 379200 446088 380000 446208 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 325048 800 325168 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 65062 479200 65118 480000 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 379200 397128 380000 397248 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 251822 479200 251878 480000 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 0 409368 800 409488 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 298834 479200 298890 480000 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 320730 479200 320786 480000 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 323306 479200 323362 480000 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 249890 0 249946 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 182914 479200 182970 480000 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 373538 0 373594 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 182928 800 183048 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 379200 132608 380000 132728 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 231888 800 232008 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 307368 800 307488 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 0 420928 800 421048 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 191088 800 191208 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 171966 479200 172022 480000 6 la_oenb[74]
port 473 nsew signal input
rlabel metal3 s 379200 4768 380000 4888 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 0 357008 800 357128 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 379200 347488 380000 347608 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 379200 440648 380000 440768 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 258408 800 258528 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 313488 800 313608 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 379200 95208 380000 95328 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 379200 417528 380000 417648 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 114006 479200 114062 480000 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 379200 356328 380000 356448 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 360014 0 360070 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 223048 800 223168 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 379200 147568 380000 147688 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 81162 479200 81218 480000 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 379200 59848 380000 59968 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 0 397808 800 397928 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 167968 800 168088 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 263414 0 263470 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 379200 414128 380000 414248 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 379200 65968 380000 66088 6 la_oenb[95]
port 496 nsew signal input
rlabel metal3 s 0 432488 800 432608 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 218978 479200 219034 480000 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 0 417528 800 417648 6 la_oenb[99]
port 500 nsew signal input
rlabel metal3 s 0 461048 800 461168 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 477680 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 477680 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 477680 6 vssd1
port 503 nsew ground input
rlabel metal3 s 379200 173408 380000 173528 6 wb_clk_i
port 504 nsew signal input
rlabel metal3 s 0 391688 800 391808 6 wb_rst_i
port 505 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 139122 479200 139178 480000 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 42522 479200 42578 480000 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal3 s 0 336608 800 336728 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal3 s 0 261128 800 261248 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal3 s 379200 437928 380000 438048 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal3 s 379200 408688 380000 408808 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 291106 0 291162 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal3 s 379200 231208 380000 231328 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal3 s 379200 63248 380000 63368 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 144274 479200 144330 480000 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 273718 479200 273774 480000 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 258262 0 258318 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 368386 0 368442 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal3 s 379200 187688 380000 187808 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal3 s 0 388968 800 389088 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 15474 479200 15530 480000 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal3 s 379200 350208 380000 350328 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 334254 479200 334310 480000 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 224130 479200 224186 480000 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal3 s 379200 272008 380000 272128 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 349066 0 349122 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 215758 479200 215814 480000 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 334898 0 334954 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal3 s 379200 68688 380000 68808 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal3 s 379200 196528 380000 196648 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 20626 479200 20682 480000 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal3 s 379200 478048 380000 478168 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal3 s 0 252288 800 252408 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal3 s 0 286968 800 287088 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal3 s 379200 310088 380000 310208 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 193862 479200 193918 480000 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 301410 479200 301466 480000 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal3 s 0 394408 800 394528 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal3 s 379200 342048 380000 342168 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 317510 479200 317566 480000 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal3 s 0 188368 800 188488 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal3 s 379200 422968 380000 423088 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal3 s 379200 211488 380000 211608 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 271142 479200 271198 480000 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 12254 479200 12310 480000 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal3 s 379200 335928 380000 336048 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 357438 0 357494 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal3 s 379200 193808 380000 193928 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal3 s 0 174088 800 174208 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal3 s 379200 74808 380000 74928 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal3 s 379200 255008 380000 255128 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 262770 479200 262826 480000 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal3 s 379200 463768 380000 463888 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal3 s 379200 77528 380000 77648 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal3 s 379200 312808 380000 312928 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal3 s 379200 469888 380000 470008 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 249246 479200 249302 480000 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal3 s 379200 104048 380000 104168 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 288530 0 288586 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 338118 0 338174 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal3 s 0 353608 800 353728 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 56690 479200 56746 480000 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 163594 479200 163650 480000 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 67638 479200 67694 480000 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 230570 0 230626 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 238298 479200 238354 480000 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal3 s 379200 170688 380000 170808 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal3 s 0 272688 800 272808 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal3 s 379200 388288 380000 388408 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal3 s 379200 370608 380000 370728 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 255686 0 255742 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 229926 479200 229982 480000 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 227350 479200 227406 480000 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal3 s 0 400528 800 400648 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 1306 479200 1362 480000 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 302054 0 302110 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal3 s 0 362448 800 362568 6 wbs_stb_i
port 608 nsew signal input
rlabel metal3 s 379200 257728 380000 257848 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 380000 480000
string LEFview TRUE
string GDS_FILE /home/shahid/caravel_user_project/openlane/user_proj_systollic/runs/user_proj_systollic/results/magic/user_proj_systollic.gds
string GDS_END 50064914
string GDS_START 501748
<< end >>

