VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OpampM
  CLASS BLOCK ;
  FOREIGN OpampM ;
  ORIGIN 46.105 50.020 ;
  SIZE 151.125 BY 107.390 ;
  PIN VN
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER li1 ;
        RECT 2.600 2.975 18.110 3.295 ;
      LAYER mcon ;
        RECT 2.855 3.055 3.025 3.225 ;
        RECT 3.215 3.055 3.385 3.225 ;
        RECT 3.575 3.055 3.745 3.225 ;
        RECT 3.935 3.055 4.105 3.225 ;
        RECT 4.295 3.055 4.465 3.225 ;
        RECT 4.655 3.055 4.825 3.225 ;
        RECT 5.015 3.055 5.185 3.225 ;
        RECT 5.375 3.055 5.545 3.225 ;
        RECT 5.735 3.055 5.905 3.225 ;
        RECT 6.095 3.055 6.265 3.225 ;
        RECT 6.455 3.055 6.625 3.225 ;
        RECT 6.815 3.055 6.985 3.225 ;
        RECT 7.175 3.055 7.345 3.225 ;
        RECT 7.535 3.055 7.705 3.225 ;
        RECT 7.895 3.055 8.065 3.225 ;
        RECT 8.255 3.055 8.425 3.225 ;
        RECT 8.615 3.055 8.785 3.225 ;
        RECT 8.975 3.055 9.145 3.225 ;
        RECT 9.335 3.055 9.505 3.225 ;
        RECT 9.695 3.055 9.865 3.225 ;
        RECT 10.055 3.055 10.225 3.225 ;
        RECT 10.415 3.055 10.585 3.225 ;
        RECT 10.775 3.055 10.945 3.225 ;
        RECT 11.135 3.055 11.305 3.225 ;
        RECT 11.495 3.055 11.665 3.225 ;
        RECT 11.855 3.055 12.025 3.225 ;
        RECT 12.215 3.055 12.385 3.225 ;
        RECT 12.575 3.055 12.745 3.225 ;
        RECT 12.935 3.055 13.105 3.225 ;
        RECT 13.295 3.055 13.465 3.225 ;
        RECT 13.655 3.055 13.825 3.225 ;
        RECT 14.015 3.055 14.185 3.225 ;
        RECT 14.375 3.055 14.545 3.225 ;
        RECT 14.735 3.055 14.905 3.225 ;
        RECT 15.095 3.055 15.265 3.225 ;
        RECT 15.455 3.055 15.625 3.225 ;
        RECT 15.815 3.055 15.985 3.225 ;
        RECT 16.175 3.055 16.345 3.225 ;
        RECT 16.535 3.055 16.705 3.225 ;
        RECT 16.895 3.055 17.065 3.225 ;
        RECT 17.255 3.055 17.425 3.225 ;
        RECT 17.615 3.055 17.785 3.225 ;
      LAYER met1 ;
        RECT -5.225 3.295 -0.720 4.680 ;
        RECT -5.225 2.975 18.110 3.295 ;
        RECT -5.225 1.205 -0.720 2.975 ;
      LAYER via ;
        RECT -4.735 1.665 -1.275 4.165 ;
      LAYER met2 ;
        RECT -46.105 1.205 -0.720 4.680 ;
    END
  END VN
  PIN VP
    ANTENNAGATEAREA 25.000000 ;
    PORT
      LAYER li1 ;
        RECT 3.390 8.975 17.320 9.295 ;
      LAYER mcon ;
        RECT 3.530 9.055 3.700 9.225 ;
        RECT 3.890 9.055 4.060 9.225 ;
        RECT 4.250 9.055 4.420 9.225 ;
        RECT 4.610 9.055 4.780 9.225 ;
        RECT 4.970 9.055 5.140 9.225 ;
        RECT 5.330 9.055 5.500 9.225 ;
        RECT 5.690 9.055 5.860 9.225 ;
        RECT 6.050 9.055 6.220 9.225 ;
        RECT 6.410 9.055 6.580 9.225 ;
        RECT 6.770 9.055 6.940 9.225 ;
        RECT 7.130 9.055 7.300 9.225 ;
        RECT 7.490 9.055 7.660 9.225 ;
        RECT 7.850 9.055 8.020 9.225 ;
        RECT 8.210 9.055 8.380 9.225 ;
        RECT 8.570 9.055 8.740 9.225 ;
        RECT 8.930 9.055 9.100 9.225 ;
        RECT 9.290 9.055 9.460 9.225 ;
        RECT 9.650 9.055 9.820 9.225 ;
        RECT 10.010 9.055 10.180 9.225 ;
        RECT 10.370 9.055 10.540 9.225 ;
        RECT 10.730 9.055 10.900 9.225 ;
        RECT 11.090 9.055 11.260 9.225 ;
        RECT 11.450 9.055 11.620 9.225 ;
        RECT 11.810 9.055 11.980 9.225 ;
        RECT 12.170 9.055 12.340 9.225 ;
        RECT 12.530 9.055 12.700 9.225 ;
        RECT 12.890 9.055 13.060 9.225 ;
        RECT 13.250 9.055 13.420 9.225 ;
        RECT 13.610 9.055 13.780 9.225 ;
        RECT 13.970 9.055 14.140 9.225 ;
        RECT 14.330 9.055 14.500 9.225 ;
        RECT 14.690 9.055 14.860 9.225 ;
        RECT 15.050 9.055 15.220 9.225 ;
        RECT 15.410 9.055 15.580 9.225 ;
        RECT 15.770 9.055 15.940 9.225 ;
        RECT 16.130 9.055 16.300 9.225 ;
        RECT 16.490 9.055 16.660 9.225 ;
        RECT 16.850 9.055 17.020 9.225 ;
      LAYER met1 ;
        RECT -2.920 9.295 -0.720 10.955 ;
        RECT -2.920 8.975 17.320 9.295 ;
        RECT -2.920 7.480 -0.720 8.975 ;
      LAYER via ;
        RECT -2.620 7.780 -1.080 10.600 ;
      LAYER met2 ;
        RECT -46.105 7.480 -0.720 10.955 ;
    END
  END VP
  PIN IBIAS
    ANTENNAGATEAREA 52.500000 ;
    ANTENNADIFFAREA 3.045000 ;
    PORT
      LAYER li1 ;
        RECT 3.460 -1.555 11.070 -1.235 ;
        RECT 7.970 -12.415 8.140 -1.875 ;
        RECT 3.460 -13.055 11.070 -12.735 ;
      LAYER mcon ;
        RECT 3.560 -1.475 3.730 -1.305 ;
        RECT 3.920 -1.475 4.090 -1.305 ;
        RECT 4.280 -1.475 4.450 -1.305 ;
        RECT 4.640 -1.475 4.810 -1.305 ;
        RECT 5.000 -1.475 5.170 -1.305 ;
        RECT 5.360 -1.475 5.530 -1.305 ;
        RECT 5.720 -1.475 5.890 -1.305 ;
        RECT 6.080 -1.475 6.250 -1.305 ;
        RECT 6.440 -1.475 6.610 -1.305 ;
        RECT 6.800 -1.475 6.970 -1.305 ;
        RECT 7.160 -1.475 7.330 -1.305 ;
        RECT 7.520 -1.475 7.690 -1.305 ;
        RECT 7.880 -1.475 8.050 -1.305 ;
        RECT 8.240 -1.475 8.410 -1.305 ;
        RECT 8.600 -1.475 8.770 -1.305 ;
        RECT 8.960 -1.475 9.130 -1.305 ;
        RECT 9.320 -1.475 9.490 -1.305 ;
        RECT 9.680 -1.475 9.850 -1.305 ;
        RECT 10.040 -1.475 10.210 -1.305 ;
        RECT 10.400 -1.475 10.570 -1.305 ;
        RECT 10.760 -1.475 10.930 -1.305 ;
        RECT 7.970 -2.190 8.140 -2.020 ;
        RECT 7.970 -2.550 8.140 -2.380 ;
        RECT 7.970 -2.910 8.140 -2.740 ;
        RECT 7.970 -3.270 8.140 -3.100 ;
        RECT 7.970 -3.630 8.140 -3.460 ;
        RECT 7.970 -3.990 8.140 -3.820 ;
        RECT 7.970 -4.350 8.140 -4.180 ;
        RECT 7.970 -4.710 8.140 -4.540 ;
        RECT 7.970 -5.070 8.140 -4.900 ;
        RECT 7.970 -5.430 8.140 -5.260 ;
        RECT 7.970 -5.790 8.140 -5.620 ;
        RECT 7.970 -6.150 8.140 -5.980 ;
        RECT 7.970 -6.510 8.140 -6.340 ;
        RECT 7.970 -6.870 8.140 -6.700 ;
        RECT 7.970 -7.230 8.140 -7.060 ;
        RECT 7.970 -7.590 8.140 -7.420 ;
        RECT 7.970 -7.950 8.140 -7.780 ;
        RECT 7.970 -8.310 8.140 -8.140 ;
        RECT 7.970 -8.670 8.140 -8.500 ;
        RECT 7.970 -9.030 8.140 -8.860 ;
        RECT 7.970 -9.390 8.140 -9.220 ;
        RECT 7.970 -9.750 8.140 -9.580 ;
        RECT 7.970 -10.110 8.140 -9.940 ;
        RECT 7.970 -10.470 8.140 -10.300 ;
        RECT 7.970 -10.830 8.140 -10.660 ;
        RECT 7.970 -11.190 8.140 -11.020 ;
        RECT 7.970 -11.550 8.140 -11.380 ;
        RECT 7.970 -11.910 8.140 -11.740 ;
        RECT 7.970 -12.270 8.140 -12.100 ;
        RECT 3.560 -12.975 3.730 -12.805 ;
        RECT 3.920 -12.975 4.090 -12.805 ;
        RECT 4.280 -12.975 4.450 -12.805 ;
        RECT 4.640 -12.975 4.810 -12.805 ;
        RECT 5.000 -12.975 5.170 -12.805 ;
        RECT 5.360 -12.975 5.530 -12.805 ;
        RECT 5.720 -12.975 5.890 -12.805 ;
        RECT 6.080 -12.975 6.250 -12.805 ;
        RECT 6.440 -12.975 6.610 -12.805 ;
        RECT 6.800 -12.975 6.970 -12.805 ;
        RECT 7.160 -12.975 7.330 -12.805 ;
        RECT 7.520 -12.975 7.690 -12.805 ;
        RECT 7.880 -12.975 8.050 -12.805 ;
        RECT 8.240 -12.975 8.410 -12.805 ;
        RECT 8.600 -12.975 8.770 -12.805 ;
        RECT 8.960 -12.975 9.130 -12.805 ;
        RECT 9.320 -12.975 9.490 -12.805 ;
        RECT 9.680 -12.975 9.850 -12.805 ;
        RECT 10.040 -12.975 10.210 -12.805 ;
        RECT 10.400 -12.975 10.570 -12.805 ;
        RECT 10.760 -12.975 10.930 -12.805 ;
      LAYER met1 ;
        RECT 2.400 -1.555 12.100 -1.235 ;
        RECT 2.400 -12.735 2.860 -1.555 ;
        RECT 7.940 -2.010 8.170 -1.895 ;
        RECT 7.895 -2.825 8.215 -2.010 ;
        RECT 7.940 -12.395 8.170 -2.825 ;
        RECT 11.640 -12.735 12.100 -1.555 ;
        RECT 2.400 -13.055 12.100 -12.735 ;
      LAYER via ;
        RECT 2.500 -2.380 2.760 -2.120 ;
        RECT 2.500 -2.700 2.760 -2.440 ;
        RECT 7.925 -2.390 8.185 -2.130 ;
        RECT 7.925 -2.710 8.185 -2.450 ;
        RECT 11.730 -2.420 11.990 -2.160 ;
        RECT 11.730 -2.740 11.990 -2.480 ;
      LAYER met2 ;
        RECT -45.880 -2.005 -0.625 -0.815 ;
        RECT -45.880 -2.835 12.100 -2.005 ;
        RECT -45.880 -4.290 -0.625 -2.835 ;
    END
  END IBIAS
  PIN VDD
    ANTENNADIFFAREA 269.293793 ;
    PORT
      LAYER nwell ;
        RECT -0.090 12.555 21.295 24.005 ;
        RECT 23.240 1.040 53.600 23.910 ;
      LAYER li1 ;
        RECT 2.680 23.650 51.925 25.620 ;
        RECT 0.715 23.400 51.925 23.650 ;
        RECT 0.715 22.745 52.255 23.400 ;
        RECT 0.715 14.340 1.805 22.745 ;
        RECT 19.515 21.720 52.255 22.745 ;
        RECT 3.480 15.550 3.650 21.590 ;
        RECT 5.060 15.550 5.230 21.590 ;
        RECT 6.640 15.550 6.810 21.590 ;
        RECT 8.220 15.550 8.390 21.590 ;
        RECT 9.800 15.550 9.970 21.590 ;
        RECT 11.380 15.550 11.550 21.590 ;
        RECT 12.960 15.550 13.130 21.590 ;
        RECT 14.540 15.550 14.710 21.590 ;
        RECT 16.120 15.550 16.290 21.590 ;
        RECT 17.700 15.550 17.870 21.590 ;
        RECT 19.515 14.340 25.565 21.720 ;
        RECT 0.715 13.435 25.565 14.340 ;
        RECT 24.145 4.260 25.565 13.435 ;
        RECT 28.265 5.725 28.435 19.965 ;
        RECT 29.845 5.725 30.015 19.965 ;
        RECT 31.425 5.725 31.595 19.965 ;
        RECT 33.005 5.725 33.175 19.965 ;
        RECT 34.585 5.725 34.755 19.965 ;
        RECT 36.165 5.725 36.335 19.965 ;
        RECT 37.745 5.725 37.915 19.965 ;
        RECT 39.325 5.725 39.495 19.965 ;
        RECT 40.905 5.725 41.075 19.965 ;
        RECT 42.485 5.725 42.655 19.965 ;
        RECT 44.065 5.725 44.235 19.965 ;
        RECT 45.645 5.725 45.815 19.965 ;
        RECT 47.225 5.725 47.395 19.965 ;
        RECT 50.835 4.260 52.255 21.720 ;
        RECT 24.145 2.580 52.255 4.260 ;
      LAYER mcon ;
        RECT 2.885 22.845 51.655 25.535 ;
        RECT 0.805 18.375 0.975 18.545 ;
        RECT 1.165 18.375 1.335 18.545 ;
        RECT 1.525 18.375 1.695 18.545 ;
        RECT 3.480 21.185 3.650 21.355 ;
        RECT 3.480 20.825 3.650 20.995 ;
        RECT 3.480 20.465 3.650 20.635 ;
        RECT 3.480 20.105 3.650 20.275 ;
        RECT 3.480 19.745 3.650 19.915 ;
        RECT 3.480 19.385 3.650 19.555 ;
        RECT 3.480 19.025 3.650 19.195 ;
        RECT 3.480 18.665 3.650 18.835 ;
        RECT 3.480 18.305 3.650 18.475 ;
        RECT 3.480 17.945 3.650 18.115 ;
        RECT 3.480 17.585 3.650 17.755 ;
        RECT 3.480 17.225 3.650 17.395 ;
        RECT 3.480 16.865 3.650 17.035 ;
        RECT 3.480 16.505 3.650 16.675 ;
        RECT 3.480 16.145 3.650 16.315 ;
        RECT 3.480 15.785 3.650 15.955 ;
        RECT 5.060 21.185 5.230 21.355 ;
        RECT 5.060 20.825 5.230 20.995 ;
        RECT 5.060 20.465 5.230 20.635 ;
        RECT 5.060 20.105 5.230 20.275 ;
        RECT 5.060 19.745 5.230 19.915 ;
        RECT 5.060 19.385 5.230 19.555 ;
        RECT 5.060 19.025 5.230 19.195 ;
        RECT 5.060 18.665 5.230 18.835 ;
        RECT 5.060 18.305 5.230 18.475 ;
        RECT 5.060 17.945 5.230 18.115 ;
        RECT 5.060 17.585 5.230 17.755 ;
        RECT 5.060 17.225 5.230 17.395 ;
        RECT 5.060 16.865 5.230 17.035 ;
        RECT 5.060 16.505 5.230 16.675 ;
        RECT 5.060 16.145 5.230 16.315 ;
        RECT 5.060 15.785 5.230 15.955 ;
        RECT 6.640 21.185 6.810 21.355 ;
        RECT 6.640 20.825 6.810 20.995 ;
        RECT 6.640 20.465 6.810 20.635 ;
        RECT 6.640 20.105 6.810 20.275 ;
        RECT 6.640 19.745 6.810 19.915 ;
        RECT 6.640 19.385 6.810 19.555 ;
        RECT 6.640 19.025 6.810 19.195 ;
        RECT 6.640 18.665 6.810 18.835 ;
        RECT 6.640 18.305 6.810 18.475 ;
        RECT 6.640 17.945 6.810 18.115 ;
        RECT 6.640 17.585 6.810 17.755 ;
        RECT 6.640 17.225 6.810 17.395 ;
        RECT 6.640 16.865 6.810 17.035 ;
        RECT 6.640 16.505 6.810 16.675 ;
        RECT 6.640 16.145 6.810 16.315 ;
        RECT 6.640 15.785 6.810 15.955 ;
        RECT 8.220 21.185 8.390 21.355 ;
        RECT 8.220 20.825 8.390 20.995 ;
        RECT 8.220 20.465 8.390 20.635 ;
        RECT 8.220 20.105 8.390 20.275 ;
        RECT 8.220 19.745 8.390 19.915 ;
        RECT 8.220 19.385 8.390 19.555 ;
        RECT 8.220 19.025 8.390 19.195 ;
        RECT 8.220 18.665 8.390 18.835 ;
        RECT 8.220 18.305 8.390 18.475 ;
        RECT 8.220 17.945 8.390 18.115 ;
        RECT 8.220 17.585 8.390 17.755 ;
        RECT 8.220 17.225 8.390 17.395 ;
        RECT 8.220 16.865 8.390 17.035 ;
        RECT 8.220 16.505 8.390 16.675 ;
        RECT 8.220 16.145 8.390 16.315 ;
        RECT 8.220 15.785 8.390 15.955 ;
        RECT 9.800 21.185 9.970 21.355 ;
        RECT 9.800 20.825 9.970 20.995 ;
        RECT 9.800 20.465 9.970 20.635 ;
        RECT 9.800 20.105 9.970 20.275 ;
        RECT 9.800 19.745 9.970 19.915 ;
        RECT 9.800 19.385 9.970 19.555 ;
        RECT 9.800 19.025 9.970 19.195 ;
        RECT 9.800 18.665 9.970 18.835 ;
        RECT 9.800 18.305 9.970 18.475 ;
        RECT 9.800 17.945 9.970 18.115 ;
        RECT 9.800 17.585 9.970 17.755 ;
        RECT 9.800 17.225 9.970 17.395 ;
        RECT 9.800 16.865 9.970 17.035 ;
        RECT 9.800 16.505 9.970 16.675 ;
        RECT 9.800 16.145 9.970 16.315 ;
        RECT 9.800 15.785 9.970 15.955 ;
        RECT 11.380 21.185 11.550 21.355 ;
        RECT 11.380 20.825 11.550 20.995 ;
        RECT 11.380 20.465 11.550 20.635 ;
        RECT 11.380 20.105 11.550 20.275 ;
        RECT 11.380 19.745 11.550 19.915 ;
        RECT 11.380 19.385 11.550 19.555 ;
        RECT 11.380 19.025 11.550 19.195 ;
        RECT 11.380 18.665 11.550 18.835 ;
        RECT 11.380 18.305 11.550 18.475 ;
        RECT 11.380 17.945 11.550 18.115 ;
        RECT 11.380 17.585 11.550 17.755 ;
        RECT 11.380 17.225 11.550 17.395 ;
        RECT 11.380 16.865 11.550 17.035 ;
        RECT 11.380 16.505 11.550 16.675 ;
        RECT 11.380 16.145 11.550 16.315 ;
        RECT 11.380 15.785 11.550 15.955 ;
        RECT 12.960 21.185 13.130 21.355 ;
        RECT 12.960 20.825 13.130 20.995 ;
        RECT 12.960 20.465 13.130 20.635 ;
        RECT 12.960 20.105 13.130 20.275 ;
        RECT 12.960 19.745 13.130 19.915 ;
        RECT 12.960 19.385 13.130 19.555 ;
        RECT 12.960 19.025 13.130 19.195 ;
        RECT 12.960 18.665 13.130 18.835 ;
        RECT 12.960 18.305 13.130 18.475 ;
        RECT 12.960 17.945 13.130 18.115 ;
        RECT 12.960 17.585 13.130 17.755 ;
        RECT 12.960 17.225 13.130 17.395 ;
        RECT 12.960 16.865 13.130 17.035 ;
        RECT 12.960 16.505 13.130 16.675 ;
        RECT 12.960 16.145 13.130 16.315 ;
        RECT 12.960 15.785 13.130 15.955 ;
        RECT 14.540 21.185 14.710 21.355 ;
        RECT 14.540 20.825 14.710 20.995 ;
        RECT 14.540 20.465 14.710 20.635 ;
        RECT 14.540 20.105 14.710 20.275 ;
        RECT 14.540 19.745 14.710 19.915 ;
        RECT 14.540 19.385 14.710 19.555 ;
        RECT 14.540 19.025 14.710 19.195 ;
        RECT 14.540 18.665 14.710 18.835 ;
        RECT 14.540 18.305 14.710 18.475 ;
        RECT 14.540 17.945 14.710 18.115 ;
        RECT 14.540 17.585 14.710 17.755 ;
        RECT 14.540 17.225 14.710 17.395 ;
        RECT 14.540 16.865 14.710 17.035 ;
        RECT 14.540 16.505 14.710 16.675 ;
        RECT 14.540 16.145 14.710 16.315 ;
        RECT 14.540 15.785 14.710 15.955 ;
        RECT 16.120 21.185 16.290 21.355 ;
        RECT 16.120 20.825 16.290 20.995 ;
        RECT 16.120 20.465 16.290 20.635 ;
        RECT 16.120 20.105 16.290 20.275 ;
        RECT 16.120 19.745 16.290 19.915 ;
        RECT 16.120 19.385 16.290 19.555 ;
        RECT 16.120 19.025 16.290 19.195 ;
        RECT 16.120 18.665 16.290 18.835 ;
        RECT 16.120 18.305 16.290 18.475 ;
        RECT 16.120 17.945 16.290 18.115 ;
        RECT 16.120 17.585 16.290 17.755 ;
        RECT 16.120 17.225 16.290 17.395 ;
        RECT 16.120 16.865 16.290 17.035 ;
        RECT 16.120 16.505 16.290 16.675 ;
        RECT 16.120 16.145 16.290 16.315 ;
        RECT 16.120 15.785 16.290 15.955 ;
        RECT 17.700 21.185 17.870 21.355 ;
        RECT 17.700 20.825 17.870 20.995 ;
        RECT 17.700 20.465 17.870 20.635 ;
        RECT 17.700 20.105 17.870 20.275 ;
        RECT 17.700 19.745 17.870 19.915 ;
        RECT 17.700 19.385 17.870 19.555 ;
        RECT 17.700 19.025 17.870 19.195 ;
        RECT 17.700 18.665 17.870 18.835 ;
        RECT 17.700 18.305 17.870 18.475 ;
        RECT 17.700 17.945 17.870 18.115 ;
        RECT 17.700 17.585 17.870 17.755 ;
        RECT 17.700 17.225 17.870 17.395 ;
        RECT 17.700 16.865 17.870 17.035 ;
        RECT 17.700 16.505 17.870 16.675 ;
        RECT 17.700 16.145 17.870 16.315 ;
        RECT 17.700 15.785 17.870 15.955 ;
        RECT 19.610 18.380 19.780 18.550 ;
        RECT 19.970 18.380 20.140 18.550 ;
        RECT 20.330 18.380 20.500 18.550 ;
        RECT 24.420 16.325 25.310 19.375 ;
        RECT 28.265 19.600 28.435 19.770 ;
        RECT 28.265 19.240 28.435 19.410 ;
        RECT 28.265 18.880 28.435 19.050 ;
        RECT 28.265 18.520 28.435 18.690 ;
        RECT 28.265 18.160 28.435 18.330 ;
        RECT 28.265 17.800 28.435 17.970 ;
        RECT 28.265 17.440 28.435 17.610 ;
        RECT 28.265 17.080 28.435 17.250 ;
        RECT 28.265 16.720 28.435 16.890 ;
        RECT 28.265 16.360 28.435 16.530 ;
        RECT 28.265 16.000 28.435 16.170 ;
        RECT 28.265 15.640 28.435 15.810 ;
        RECT 28.265 15.280 28.435 15.450 ;
        RECT 28.265 14.920 28.435 15.090 ;
        RECT 28.265 14.560 28.435 14.730 ;
        RECT 28.265 14.200 28.435 14.370 ;
        RECT 28.265 13.840 28.435 14.010 ;
        RECT 28.265 13.480 28.435 13.650 ;
        RECT 28.265 13.120 28.435 13.290 ;
        RECT 28.265 12.760 28.435 12.930 ;
        RECT 28.265 12.400 28.435 12.570 ;
        RECT 28.265 12.040 28.435 12.210 ;
        RECT 28.265 11.680 28.435 11.850 ;
        RECT 28.265 11.320 28.435 11.490 ;
        RECT 28.265 10.960 28.435 11.130 ;
        RECT 28.265 10.600 28.435 10.770 ;
        RECT 28.265 10.240 28.435 10.410 ;
        RECT 28.265 9.880 28.435 10.050 ;
        RECT 28.265 9.520 28.435 9.690 ;
        RECT 28.265 9.160 28.435 9.330 ;
        RECT 28.265 8.800 28.435 8.970 ;
        RECT 28.265 8.440 28.435 8.610 ;
        RECT 28.265 8.080 28.435 8.250 ;
        RECT 28.265 7.720 28.435 7.890 ;
        RECT 28.265 7.360 28.435 7.530 ;
        RECT 28.265 7.000 28.435 7.170 ;
        RECT 28.265 6.640 28.435 6.810 ;
        RECT 28.265 6.280 28.435 6.450 ;
        RECT 28.265 5.920 28.435 6.090 ;
        RECT 29.845 19.600 30.015 19.770 ;
        RECT 29.845 19.240 30.015 19.410 ;
        RECT 29.845 18.880 30.015 19.050 ;
        RECT 29.845 18.520 30.015 18.690 ;
        RECT 29.845 18.160 30.015 18.330 ;
        RECT 29.845 17.800 30.015 17.970 ;
        RECT 29.845 17.440 30.015 17.610 ;
        RECT 29.845 17.080 30.015 17.250 ;
        RECT 29.845 16.720 30.015 16.890 ;
        RECT 29.845 16.360 30.015 16.530 ;
        RECT 29.845 16.000 30.015 16.170 ;
        RECT 29.845 15.640 30.015 15.810 ;
        RECT 29.845 15.280 30.015 15.450 ;
        RECT 29.845 14.920 30.015 15.090 ;
        RECT 29.845 14.560 30.015 14.730 ;
        RECT 29.845 14.200 30.015 14.370 ;
        RECT 29.845 13.840 30.015 14.010 ;
        RECT 29.845 13.480 30.015 13.650 ;
        RECT 29.845 13.120 30.015 13.290 ;
        RECT 29.845 12.760 30.015 12.930 ;
        RECT 29.845 12.400 30.015 12.570 ;
        RECT 29.845 12.040 30.015 12.210 ;
        RECT 29.845 11.680 30.015 11.850 ;
        RECT 29.845 11.320 30.015 11.490 ;
        RECT 29.845 10.960 30.015 11.130 ;
        RECT 29.845 10.600 30.015 10.770 ;
        RECT 29.845 10.240 30.015 10.410 ;
        RECT 29.845 9.880 30.015 10.050 ;
        RECT 29.845 9.520 30.015 9.690 ;
        RECT 29.845 9.160 30.015 9.330 ;
        RECT 29.845 8.800 30.015 8.970 ;
        RECT 29.845 8.440 30.015 8.610 ;
        RECT 29.845 8.080 30.015 8.250 ;
        RECT 29.845 7.720 30.015 7.890 ;
        RECT 29.845 7.360 30.015 7.530 ;
        RECT 29.845 7.000 30.015 7.170 ;
        RECT 29.845 6.640 30.015 6.810 ;
        RECT 29.845 6.280 30.015 6.450 ;
        RECT 29.845 5.920 30.015 6.090 ;
        RECT 31.425 19.600 31.595 19.770 ;
        RECT 31.425 19.240 31.595 19.410 ;
        RECT 31.425 18.880 31.595 19.050 ;
        RECT 31.425 18.520 31.595 18.690 ;
        RECT 31.425 18.160 31.595 18.330 ;
        RECT 31.425 17.800 31.595 17.970 ;
        RECT 31.425 17.440 31.595 17.610 ;
        RECT 31.425 17.080 31.595 17.250 ;
        RECT 31.425 16.720 31.595 16.890 ;
        RECT 31.425 16.360 31.595 16.530 ;
        RECT 31.425 16.000 31.595 16.170 ;
        RECT 31.425 15.640 31.595 15.810 ;
        RECT 31.425 15.280 31.595 15.450 ;
        RECT 31.425 14.920 31.595 15.090 ;
        RECT 31.425 14.560 31.595 14.730 ;
        RECT 31.425 14.200 31.595 14.370 ;
        RECT 31.425 13.840 31.595 14.010 ;
        RECT 31.425 13.480 31.595 13.650 ;
        RECT 31.425 13.120 31.595 13.290 ;
        RECT 31.425 12.760 31.595 12.930 ;
        RECT 31.425 12.400 31.595 12.570 ;
        RECT 31.425 12.040 31.595 12.210 ;
        RECT 31.425 11.680 31.595 11.850 ;
        RECT 31.425 11.320 31.595 11.490 ;
        RECT 31.425 10.960 31.595 11.130 ;
        RECT 31.425 10.600 31.595 10.770 ;
        RECT 31.425 10.240 31.595 10.410 ;
        RECT 31.425 9.880 31.595 10.050 ;
        RECT 31.425 9.520 31.595 9.690 ;
        RECT 31.425 9.160 31.595 9.330 ;
        RECT 31.425 8.800 31.595 8.970 ;
        RECT 31.425 8.440 31.595 8.610 ;
        RECT 31.425 8.080 31.595 8.250 ;
        RECT 31.425 7.720 31.595 7.890 ;
        RECT 31.425 7.360 31.595 7.530 ;
        RECT 31.425 7.000 31.595 7.170 ;
        RECT 31.425 6.640 31.595 6.810 ;
        RECT 31.425 6.280 31.595 6.450 ;
        RECT 31.425 5.920 31.595 6.090 ;
        RECT 33.005 19.600 33.175 19.770 ;
        RECT 33.005 19.240 33.175 19.410 ;
        RECT 33.005 18.880 33.175 19.050 ;
        RECT 33.005 18.520 33.175 18.690 ;
        RECT 33.005 18.160 33.175 18.330 ;
        RECT 33.005 17.800 33.175 17.970 ;
        RECT 33.005 17.440 33.175 17.610 ;
        RECT 33.005 17.080 33.175 17.250 ;
        RECT 33.005 16.720 33.175 16.890 ;
        RECT 33.005 16.360 33.175 16.530 ;
        RECT 33.005 16.000 33.175 16.170 ;
        RECT 33.005 15.640 33.175 15.810 ;
        RECT 33.005 15.280 33.175 15.450 ;
        RECT 33.005 14.920 33.175 15.090 ;
        RECT 33.005 14.560 33.175 14.730 ;
        RECT 33.005 14.200 33.175 14.370 ;
        RECT 33.005 13.840 33.175 14.010 ;
        RECT 33.005 13.480 33.175 13.650 ;
        RECT 33.005 13.120 33.175 13.290 ;
        RECT 33.005 12.760 33.175 12.930 ;
        RECT 33.005 12.400 33.175 12.570 ;
        RECT 33.005 12.040 33.175 12.210 ;
        RECT 33.005 11.680 33.175 11.850 ;
        RECT 33.005 11.320 33.175 11.490 ;
        RECT 33.005 10.960 33.175 11.130 ;
        RECT 33.005 10.600 33.175 10.770 ;
        RECT 33.005 10.240 33.175 10.410 ;
        RECT 33.005 9.880 33.175 10.050 ;
        RECT 33.005 9.520 33.175 9.690 ;
        RECT 33.005 9.160 33.175 9.330 ;
        RECT 33.005 8.800 33.175 8.970 ;
        RECT 33.005 8.440 33.175 8.610 ;
        RECT 33.005 8.080 33.175 8.250 ;
        RECT 33.005 7.720 33.175 7.890 ;
        RECT 33.005 7.360 33.175 7.530 ;
        RECT 33.005 7.000 33.175 7.170 ;
        RECT 33.005 6.640 33.175 6.810 ;
        RECT 33.005 6.280 33.175 6.450 ;
        RECT 33.005 5.920 33.175 6.090 ;
        RECT 34.585 19.600 34.755 19.770 ;
        RECT 34.585 19.240 34.755 19.410 ;
        RECT 34.585 18.880 34.755 19.050 ;
        RECT 34.585 18.520 34.755 18.690 ;
        RECT 34.585 18.160 34.755 18.330 ;
        RECT 34.585 17.800 34.755 17.970 ;
        RECT 34.585 17.440 34.755 17.610 ;
        RECT 34.585 17.080 34.755 17.250 ;
        RECT 34.585 16.720 34.755 16.890 ;
        RECT 34.585 16.360 34.755 16.530 ;
        RECT 34.585 16.000 34.755 16.170 ;
        RECT 34.585 15.640 34.755 15.810 ;
        RECT 34.585 15.280 34.755 15.450 ;
        RECT 34.585 14.920 34.755 15.090 ;
        RECT 34.585 14.560 34.755 14.730 ;
        RECT 34.585 14.200 34.755 14.370 ;
        RECT 34.585 13.840 34.755 14.010 ;
        RECT 34.585 13.480 34.755 13.650 ;
        RECT 34.585 13.120 34.755 13.290 ;
        RECT 34.585 12.760 34.755 12.930 ;
        RECT 34.585 12.400 34.755 12.570 ;
        RECT 34.585 12.040 34.755 12.210 ;
        RECT 34.585 11.680 34.755 11.850 ;
        RECT 34.585 11.320 34.755 11.490 ;
        RECT 34.585 10.960 34.755 11.130 ;
        RECT 34.585 10.600 34.755 10.770 ;
        RECT 34.585 10.240 34.755 10.410 ;
        RECT 34.585 9.880 34.755 10.050 ;
        RECT 34.585 9.520 34.755 9.690 ;
        RECT 34.585 9.160 34.755 9.330 ;
        RECT 34.585 8.800 34.755 8.970 ;
        RECT 34.585 8.440 34.755 8.610 ;
        RECT 34.585 8.080 34.755 8.250 ;
        RECT 34.585 7.720 34.755 7.890 ;
        RECT 34.585 7.360 34.755 7.530 ;
        RECT 34.585 7.000 34.755 7.170 ;
        RECT 34.585 6.640 34.755 6.810 ;
        RECT 34.585 6.280 34.755 6.450 ;
        RECT 34.585 5.920 34.755 6.090 ;
        RECT 36.165 19.600 36.335 19.770 ;
        RECT 36.165 19.240 36.335 19.410 ;
        RECT 36.165 18.880 36.335 19.050 ;
        RECT 36.165 18.520 36.335 18.690 ;
        RECT 36.165 18.160 36.335 18.330 ;
        RECT 36.165 17.800 36.335 17.970 ;
        RECT 36.165 17.440 36.335 17.610 ;
        RECT 36.165 17.080 36.335 17.250 ;
        RECT 36.165 16.720 36.335 16.890 ;
        RECT 36.165 16.360 36.335 16.530 ;
        RECT 36.165 16.000 36.335 16.170 ;
        RECT 36.165 15.640 36.335 15.810 ;
        RECT 36.165 15.280 36.335 15.450 ;
        RECT 36.165 14.920 36.335 15.090 ;
        RECT 36.165 14.560 36.335 14.730 ;
        RECT 36.165 14.200 36.335 14.370 ;
        RECT 36.165 13.840 36.335 14.010 ;
        RECT 36.165 13.480 36.335 13.650 ;
        RECT 36.165 13.120 36.335 13.290 ;
        RECT 36.165 12.760 36.335 12.930 ;
        RECT 36.165 12.400 36.335 12.570 ;
        RECT 36.165 12.040 36.335 12.210 ;
        RECT 36.165 11.680 36.335 11.850 ;
        RECT 36.165 11.320 36.335 11.490 ;
        RECT 36.165 10.960 36.335 11.130 ;
        RECT 36.165 10.600 36.335 10.770 ;
        RECT 36.165 10.240 36.335 10.410 ;
        RECT 36.165 9.880 36.335 10.050 ;
        RECT 36.165 9.520 36.335 9.690 ;
        RECT 36.165 9.160 36.335 9.330 ;
        RECT 36.165 8.800 36.335 8.970 ;
        RECT 36.165 8.440 36.335 8.610 ;
        RECT 36.165 8.080 36.335 8.250 ;
        RECT 36.165 7.720 36.335 7.890 ;
        RECT 36.165 7.360 36.335 7.530 ;
        RECT 36.165 7.000 36.335 7.170 ;
        RECT 36.165 6.640 36.335 6.810 ;
        RECT 36.165 6.280 36.335 6.450 ;
        RECT 36.165 5.920 36.335 6.090 ;
        RECT 37.745 19.600 37.915 19.770 ;
        RECT 37.745 19.240 37.915 19.410 ;
        RECT 37.745 18.880 37.915 19.050 ;
        RECT 37.745 18.520 37.915 18.690 ;
        RECT 37.745 18.160 37.915 18.330 ;
        RECT 37.745 17.800 37.915 17.970 ;
        RECT 37.745 17.440 37.915 17.610 ;
        RECT 37.745 17.080 37.915 17.250 ;
        RECT 37.745 16.720 37.915 16.890 ;
        RECT 37.745 16.360 37.915 16.530 ;
        RECT 37.745 16.000 37.915 16.170 ;
        RECT 37.745 15.640 37.915 15.810 ;
        RECT 37.745 15.280 37.915 15.450 ;
        RECT 37.745 14.920 37.915 15.090 ;
        RECT 37.745 14.560 37.915 14.730 ;
        RECT 37.745 14.200 37.915 14.370 ;
        RECT 37.745 13.840 37.915 14.010 ;
        RECT 37.745 13.480 37.915 13.650 ;
        RECT 37.745 13.120 37.915 13.290 ;
        RECT 37.745 12.760 37.915 12.930 ;
        RECT 37.745 12.400 37.915 12.570 ;
        RECT 37.745 12.040 37.915 12.210 ;
        RECT 37.745 11.680 37.915 11.850 ;
        RECT 37.745 11.320 37.915 11.490 ;
        RECT 37.745 10.960 37.915 11.130 ;
        RECT 37.745 10.600 37.915 10.770 ;
        RECT 37.745 10.240 37.915 10.410 ;
        RECT 37.745 9.880 37.915 10.050 ;
        RECT 37.745 9.520 37.915 9.690 ;
        RECT 37.745 9.160 37.915 9.330 ;
        RECT 37.745 8.800 37.915 8.970 ;
        RECT 37.745 8.440 37.915 8.610 ;
        RECT 37.745 8.080 37.915 8.250 ;
        RECT 37.745 7.720 37.915 7.890 ;
        RECT 37.745 7.360 37.915 7.530 ;
        RECT 37.745 7.000 37.915 7.170 ;
        RECT 37.745 6.640 37.915 6.810 ;
        RECT 37.745 6.280 37.915 6.450 ;
        RECT 37.745 5.920 37.915 6.090 ;
        RECT 39.325 19.600 39.495 19.770 ;
        RECT 39.325 19.240 39.495 19.410 ;
        RECT 39.325 18.880 39.495 19.050 ;
        RECT 39.325 18.520 39.495 18.690 ;
        RECT 39.325 18.160 39.495 18.330 ;
        RECT 39.325 17.800 39.495 17.970 ;
        RECT 39.325 17.440 39.495 17.610 ;
        RECT 39.325 17.080 39.495 17.250 ;
        RECT 39.325 16.720 39.495 16.890 ;
        RECT 39.325 16.360 39.495 16.530 ;
        RECT 39.325 16.000 39.495 16.170 ;
        RECT 39.325 15.640 39.495 15.810 ;
        RECT 39.325 15.280 39.495 15.450 ;
        RECT 39.325 14.920 39.495 15.090 ;
        RECT 39.325 14.560 39.495 14.730 ;
        RECT 39.325 14.200 39.495 14.370 ;
        RECT 39.325 13.840 39.495 14.010 ;
        RECT 39.325 13.480 39.495 13.650 ;
        RECT 39.325 13.120 39.495 13.290 ;
        RECT 39.325 12.760 39.495 12.930 ;
        RECT 39.325 12.400 39.495 12.570 ;
        RECT 39.325 12.040 39.495 12.210 ;
        RECT 39.325 11.680 39.495 11.850 ;
        RECT 39.325 11.320 39.495 11.490 ;
        RECT 39.325 10.960 39.495 11.130 ;
        RECT 39.325 10.600 39.495 10.770 ;
        RECT 39.325 10.240 39.495 10.410 ;
        RECT 39.325 9.880 39.495 10.050 ;
        RECT 39.325 9.520 39.495 9.690 ;
        RECT 39.325 9.160 39.495 9.330 ;
        RECT 39.325 8.800 39.495 8.970 ;
        RECT 39.325 8.440 39.495 8.610 ;
        RECT 39.325 8.080 39.495 8.250 ;
        RECT 39.325 7.720 39.495 7.890 ;
        RECT 39.325 7.360 39.495 7.530 ;
        RECT 39.325 7.000 39.495 7.170 ;
        RECT 39.325 6.640 39.495 6.810 ;
        RECT 39.325 6.280 39.495 6.450 ;
        RECT 39.325 5.920 39.495 6.090 ;
        RECT 40.905 19.600 41.075 19.770 ;
        RECT 40.905 19.240 41.075 19.410 ;
        RECT 40.905 18.880 41.075 19.050 ;
        RECT 40.905 18.520 41.075 18.690 ;
        RECT 40.905 18.160 41.075 18.330 ;
        RECT 40.905 17.800 41.075 17.970 ;
        RECT 40.905 17.440 41.075 17.610 ;
        RECT 40.905 17.080 41.075 17.250 ;
        RECT 40.905 16.720 41.075 16.890 ;
        RECT 40.905 16.360 41.075 16.530 ;
        RECT 40.905 16.000 41.075 16.170 ;
        RECT 40.905 15.640 41.075 15.810 ;
        RECT 40.905 15.280 41.075 15.450 ;
        RECT 40.905 14.920 41.075 15.090 ;
        RECT 40.905 14.560 41.075 14.730 ;
        RECT 40.905 14.200 41.075 14.370 ;
        RECT 40.905 13.840 41.075 14.010 ;
        RECT 40.905 13.480 41.075 13.650 ;
        RECT 40.905 13.120 41.075 13.290 ;
        RECT 40.905 12.760 41.075 12.930 ;
        RECT 40.905 12.400 41.075 12.570 ;
        RECT 40.905 12.040 41.075 12.210 ;
        RECT 40.905 11.680 41.075 11.850 ;
        RECT 40.905 11.320 41.075 11.490 ;
        RECT 40.905 10.960 41.075 11.130 ;
        RECT 40.905 10.600 41.075 10.770 ;
        RECT 40.905 10.240 41.075 10.410 ;
        RECT 40.905 9.880 41.075 10.050 ;
        RECT 40.905 9.520 41.075 9.690 ;
        RECT 40.905 9.160 41.075 9.330 ;
        RECT 40.905 8.800 41.075 8.970 ;
        RECT 40.905 8.440 41.075 8.610 ;
        RECT 40.905 8.080 41.075 8.250 ;
        RECT 40.905 7.720 41.075 7.890 ;
        RECT 40.905 7.360 41.075 7.530 ;
        RECT 40.905 7.000 41.075 7.170 ;
        RECT 40.905 6.640 41.075 6.810 ;
        RECT 40.905 6.280 41.075 6.450 ;
        RECT 40.905 5.920 41.075 6.090 ;
        RECT 42.485 19.600 42.655 19.770 ;
        RECT 42.485 19.240 42.655 19.410 ;
        RECT 42.485 18.880 42.655 19.050 ;
        RECT 42.485 18.520 42.655 18.690 ;
        RECT 42.485 18.160 42.655 18.330 ;
        RECT 42.485 17.800 42.655 17.970 ;
        RECT 42.485 17.440 42.655 17.610 ;
        RECT 42.485 17.080 42.655 17.250 ;
        RECT 42.485 16.720 42.655 16.890 ;
        RECT 42.485 16.360 42.655 16.530 ;
        RECT 42.485 16.000 42.655 16.170 ;
        RECT 42.485 15.640 42.655 15.810 ;
        RECT 42.485 15.280 42.655 15.450 ;
        RECT 42.485 14.920 42.655 15.090 ;
        RECT 42.485 14.560 42.655 14.730 ;
        RECT 42.485 14.200 42.655 14.370 ;
        RECT 42.485 13.840 42.655 14.010 ;
        RECT 42.485 13.480 42.655 13.650 ;
        RECT 42.485 13.120 42.655 13.290 ;
        RECT 42.485 12.760 42.655 12.930 ;
        RECT 42.485 12.400 42.655 12.570 ;
        RECT 42.485 12.040 42.655 12.210 ;
        RECT 42.485 11.680 42.655 11.850 ;
        RECT 42.485 11.320 42.655 11.490 ;
        RECT 42.485 10.960 42.655 11.130 ;
        RECT 42.485 10.600 42.655 10.770 ;
        RECT 42.485 10.240 42.655 10.410 ;
        RECT 42.485 9.880 42.655 10.050 ;
        RECT 42.485 9.520 42.655 9.690 ;
        RECT 42.485 9.160 42.655 9.330 ;
        RECT 42.485 8.800 42.655 8.970 ;
        RECT 42.485 8.440 42.655 8.610 ;
        RECT 42.485 8.080 42.655 8.250 ;
        RECT 42.485 7.720 42.655 7.890 ;
        RECT 42.485 7.360 42.655 7.530 ;
        RECT 42.485 7.000 42.655 7.170 ;
        RECT 42.485 6.640 42.655 6.810 ;
        RECT 42.485 6.280 42.655 6.450 ;
        RECT 42.485 5.920 42.655 6.090 ;
        RECT 44.065 19.600 44.235 19.770 ;
        RECT 44.065 19.240 44.235 19.410 ;
        RECT 44.065 18.880 44.235 19.050 ;
        RECT 44.065 18.520 44.235 18.690 ;
        RECT 44.065 18.160 44.235 18.330 ;
        RECT 44.065 17.800 44.235 17.970 ;
        RECT 44.065 17.440 44.235 17.610 ;
        RECT 44.065 17.080 44.235 17.250 ;
        RECT 44.065 16.720 44.235 16.890 ;
        RECT 44.065 16.360 44.235 16.530 ;
        RECT 44.065 16.000 44.235 16.170 ;
        RECT 44.065 15.640 44.235 15.810 ;
        RECT 44.065 15.280 44.235 15.450 ;
        RECT 44.065 14.920 44.235 15.090 ;
        RECT 44.065 14.560 44.235 14.730 ;
        RECT 44.065 14.200 44.235 14.370 ;
        RECT 44.065 13.840 44.235 14.010 ;
        RECT 44.065 13.480 44.235 13.650 ;
        RECT 44.065 13.120 44.235 13.290 ;
        RECT 44.065 12.760 44.235 12.930 ;
        RECT 44.065 12.400 44.235 12.570 ;
        RECT 44.065 12.040 44.235 12.210 ;
        RECT 44.065 11.680 44.235 11.850 ;
        RECT 44.065 11.320 44.235 11.490 ;
        RECT 44.065 10.960 44.235 11.130 ;
        RECT 44.065 10.600 44.235 10.770 ;
        RECT 44.065 10.240 44.235 10.410 ;
        RECT 44.065 9.880 44.235 10.050 ;
        RECT 44.065 9.520 44.235 9.690 ;
        RECT 44.065 9.160 44.235 9.330 ;
        RECT 44.065 8.800 44.235 8.970 ;
        RECT 44.065 8.440 44.235 8.610 ;
        RECT 44.065 8.080 44.235 8.250 ;
        RECT 44.065 7.720 44.235 7.890 ;
        RECT 44.065 7.360 44.235 7.530 ;
        RECT 44.065 7.000 44.235 7.170 ;
        RECT 44.065 6.640 44.235 6.810 ;
        RECT 44.065 6.280 44.235 6.450 ;
        RECT 44.065 5.920 44.235 6.090 ;
        RECT 45.645 19.600 45.815 19.770 ;
        RECT 45.645 19.240 45.815 19.410 ;
        RECT 45.645 18.880 45.815 19.050 ;
        RECT 45.645 18.520 45.815 18.690 ;
        RECT 45.645 18.160 45.815 18.330 ;
        RECT 45.645 17.800 45.815 17.970 ;
        RECT 45.645 17.440 45.815 17.610 ;
        RECT 45.645 17.080 45.815 17.250 ;
        RECT 45.645 16.720 45.815 16.890 ;
        RECT 45.645 16.360 45.815 16.530 ;
        RECT 45.645 16.000 45.815 16.170 ;
        RECT 45.645 15.640 45.815 15.810 ;
        RECT 45.645 15.280 45.815 15.450 ;
        RECT 45.645 14.920 45.815 15.090 ;
        RECT 45.645 14.560 45.815 14.730 ;
        RECT 45.645 14.200 45.815 14.370 ;
        RECT 45.645 13.840 45.815 14.010 ;
        RECT 45.645 13.480 45.815 13.650 ;
        RECT 45.645 13.120 45.815 13.290 ;
        RECT 45.645 12.760 45.815 12.930 ;
        RECT 45.645 12.400 45.815 12.570 ;
        RECT 45.645 12.040 45.815 12.210 ;
        RECT 45.645 11.680 45.815 11.850 ;
        RECT 45.645 11.320 45.815 11.490 ;
        RECT 45.645 10.960 45.815 11.130 ;
        RECT 45.645 10.600 45.815 10.770 ;
        RECT 45.645 10.240 45.815 10.410 ;
        RECT 45.645 9.880 45.815 10.050 ;
        RECT 45.645 9.520 45.815 9.690 ;
        RECT 45.645 9.160 45.815 9.330 ;
        RECT 45.645 8.800 45.815 8.970 ;
        RECT 45.645 8.440 45.815 8.610 ;
        RECT 45.645 8.080 45.815 8.250 ;
        RECT 45.645 7.720 45.815 7.890 ;
        RECT 45.645 7.360 45.815 7.530 ;
        RECT 45.645 7.000 45.815 7.170 ;
        RECT 45.645 6.640 45.815 6.810 ;
        RECT 45.645 6.280 45.815 6.450 ;
        RECT 45.645 5.920 45.815 6.090 ;
        RECT 47.225 19.600 47.395 19.770 ;
        RECT 47.225 19.240 47.395 19.410 ;
        RECT 47.225 18.880 47.395 19.050 ;
        RECT 47.225 18.520 47.395 18.690 ;
        RECT 47.225 18.160 47.395 18.330 ;
        RECT 47.225 17.800 47.395 17.970 ;
        RECT 47.225 17.440 47.395 17.610 ;
        RECT 47.225 17.080 47.395 17.250 ;
        RECT 47.225 16.720 47.395 16.890 ;
        RECT 47.225 16.360 47.395 16.530 ;
        RECT 47.225 16.000 47.395 16.170 ;
        RECT 47.225 15.640 47.395 15.810 ;
        RECT 47.225 15.280 47.395 15.450 ;
        RECT 47.225 14.920 47.395 15.090 ;
        RECT 47.225 14.560 47.395 14.730 ;
        RECT 47.225 14.200 47.395 14.370 ;
        RECT 47.225 13.840 47.395 14.010 ;
        RECT 47.225 13.480 47.395 13.650 ;
        RECT 47.225 13.120 47.395 13.290 ;
        RECT 47.225 12.760 47.395 12.930 ;
        RECT 47.225 12.400 47.395 12.570 ;
        RECT 47.225 12.040 47.395 12.210 ;
        RECT 47.225 11.680 47.395 11.850 ;
        RECT 47.225 11.320 47.395 11.490 ;
        RECT 47.225 10.960 47.395 11.130 ;
        RECT 47.225 10.600 47.395 10.770 ;
        RECT 47.225 10.240 47.395 10.410 ;
        RECT 47.225 9.880 47.395 10.050 ;
        RECT 47.225 9.520 47.395 9.690 ;
        RECT 47.225 9.160 47.395 9.330 ;
        RECT 47.225 8.800 47.395 8.970 ;
        RECT 47.225 8.440 47.395 8.610 ;
        RECT 47.225 8.080 47.395 8.250 ;
        RECT 47.225 7.720 47.395 7.890 ;
        RECT 47.225 7.360 47.395 7.530 ;
        RECT 47.225 7.000 47.395 7.170 ;
        RECT 47.225 6.640 47.395 6.810 ;
        RECT 47.225 6.280 47.395 6.450 ;
        RECT 47.225 5.920 47.395 6.090 ;
        RECT 51.105 16.380 51.995 19.430 ;
      LAYER met1 ;
        RECT 2.680 22.745 51.925 25.620 ;
        RECT 3.450 18.750 3.680 21.570 ;
        RECT 5.030 18.750 5.260 21.570 ;
        RECT 6.610 18.750 6.840 21.570 ;
        RECT 8.190 18.750 8.420 21.570 ;
        RECT 9.770 18.750 10.000 21.570 ;
        RECT 11.350 18.750 11.580 21.570 ;
        RECT 12.930 18.750 13.160 21.570 ;
        RECT 14.510 18.750 14.740 21.570 ;
        RECT 16.090 18.750 16.320 21.570 ;
        RECT 17.670 18.750 17.900 21.570 ;
        RECT 0.715 18.170 1.805 18.750 ;
        RECT 3.405 18.170 3.725 18.750 ;
        RECT 4.985 18.170 5.305 18.750 ;
        RECT 6.565 18.170 6.885 18.750 ;
        RECT 8.145 18.170 8.465 18.750 ;
        RECT 9.725 18.170 10.045 18.750 ;
        RECT 11.305 18.170 11.625 18.750 ;
        RECT 12.885 18.170 13.205 18.750 ;
        RECT 14.465 18.170 14.785 18.750 ;
        RECT 16.045 18.170 16.365 18.750 ;
        RECT 17.625 18.170 17.945 18.750 ;
        RECT 19.515 18.170 20.605 18.750 ;
        RECT 3.450 15.570 3.680 18.170 ;
        RECT 5.030 15.570 5.260 18.170 ;
        RECT 6.610 15.570 6.840 18.170 ;
        RECT 8.190 15.570 8.420 18.170 ;
        RECT 9.770 15.570 10.000 18.170 ;
        RECT 11.350 15.570 11.580 18.170 ;
        RECT 12.930 15.570 13.160 18.170 ;
        RECT 14.510 15.570 14.740 18.170 ;
        RECT 16.090 15.570 16.320 18.170 ;
        RECT 17.670 15.570 17.900 18.170 ;
        RECT 24.145 16.030 25.565 19.795 ;
        RECT 28.235 19.780 28.465 19.945 ;
        RECT 29.815 19.780 30.045 19.945 ;
        RECT 31.395 19.780 31.625 19.945 ;
        RECT 32.975 19.780 33.205 19.945 ;
        RECT 34.555 19.780 34.785 19.945 ;
        RECT 36.135 19.780 36.365 19.945 ;
        RECT 37.715 19.780 37.945 19.945 ;
        RECT 39.295 19.780 39.525 19.945 ;
        RECT 40.875 19.780 41.105 19.945 ;
        RECT 42.455 19.780 42.685 19.945 ;
        RECT 44.035 19.780 44.265 19.945 ;
        RECT 45.615 19.780 45.845 19.945 ;
        RECT 47.195 19.780 47.425 19.945 ;
        RECT 28.190 16.045 28.510 19.780 ;
        RECT 29.770 16.045 30.090 19.780 ;
        RECT 31.350 16.045 31.670 19.780 ;
        RECT 32.930 16.045 33.250 19.780 ;
        RECT 34.510 16.045 34.830 19.780 ;
        RECT 36.090 16.045 36.410 19.780 ;
        RECT 37.670 16.045 37.990 19.780 ;
        RECT 39.250 16.045 39.570 19.780 ;
        RECT 40.830 16.045 41.150 19.780 ;
        RECT 42.410 16.045 42.730 19.780 ;
        RECT 43.990 16.045 44.310 19.780 ;
        RECT 45.570 16.045 45.890 19.780 ;
        RECT 47.150 16.045 47.470 19.780 ;
        RECT 28.235 5.745 28.465 16.045 ;
        RECT 29.815 5.745 30.045 16.045 ;
        RECT 31.395 5.745 31.625 16.045 ;
        RECT 32.975 5.745 33.205 16.045 ;
        RECT 34.555 5.745 34.785 16.045 ;
        RECT 36.135 5.745 36.365 16.045 ;
        RECT 37.715 5.745 37.945 16.045 ;
        RECT 39.295 5.745 39.525 16.045 ;
        RECT 40.875 5.745 41.105 16.045 ;
        RECT 42.455 5.745 42.685 16.045 ;
        RECT 44.035 5.745 44.265 16.045 ;
        RECT 45.615 5.745 45.845 16.045 ;
        RECT 47.195 5.745 47.425 16.045 ;
        RECT 50.835 16.030 52.255 19.795 ;
      LAYER via ;
        RECT 2.820 22.940 51.720 25.440 ;
        RECT 0.800 18.330 1.060 18.590 ;
        RECT 1.120 18.330 1.380 18.590 ;
        RECT 1.440 18.330 1.700 18.590 ;
        RECT 3.435 18.330 3.695 18.590 ;
        RECT 5.015 18.330 5.275 18.590 ;
        RECT 6.595 18.330 6.855 18.590 ;
        RECT 8.175 18.330 8.435 18.590 ;
        RECT 9.755 18.330 10.015 18.590 ;
        RECT 11.335 18.330 11.595 18.590 ;
        RECT 12.915 18.330 13.175 18.590 ;
        RECT 14.495 18.330 14.755 18.590 ;
        RECT 16.075 18.330 16.335 18.590 ;
        RECT 17.655 18.330 17.915 18.590 ;
        RECT 19.605 18.335 19.865 18.595 ;
        RECT 19.925 18.335 20.185 18.595 ;
        RECT 20.245 18.335 20.505 18.595 ;
        RECT 24.415 16.280 25.315 19.420 ;
        RECT 28.220 19.380 28.480 19.640 ;
        RECT 28.220 19.060 28.480 19.320 ;
        RECT 28.220 18.740 28.480 19.000 ;
        RECT 28.220 18.420 28.480 18.680 ;
        RECT 28.220 18.100 28.480 18.360 ;
        RECT 28.220 17.780 28.480 18.040 ;
        RECT 28.220 17.460 28.480 17.720 ;
        RECT 28.220 17.140 28.480 17.400 ;
        RECT 28.220 16.820 28.480 17.080 ;
        RECT 28.220 16.500 28.480 16.760 ;
        RECT 28.220 16.180 28.480 16.440 ;
        RECT 29.800 19.380 30.060 19.640 ;
        RECT 29.800 19.060 30.060 19.320 ;
        RECT 29.800 18.740 30.060 19.000 ;
        RECT 29.800 18.420 30.060 18.680 ;
        RECT 29.800 18.100 30.060 18.360 ;
        RECT 29.800 17.780 30.060 18.040 ;
        RECT 29.800 17.460 30.060 17.720 ;
        RECT 29.800 17.140 30.060 17.400 ;
        RECT 29.800 16.820 30.060 17.080 ;
        RECT 29.800 16.500 30.060 16.760 ;
        RECT 29.800 16.180 30.060 16.440 ;
        RECT 31.380 19.380 31.640 19.640 ;
        RECT 31.380 19.060 31.640 19.320 ;
        RECT 31.380 18.740 31.640 19.000 ;
        RECT 31.380 18.420 31.640 18.680 ;
        RECT 31.380 18.100 31.640 18.360 ;
        RECT 31.380 17.780 31.640 18.040 ;
        RECT 31.380 17.460 31.640 17.720 ;
        RECT 31.380 17.140 31.640 17.400 ;
        RECT 31.380 16.820 31.640 17.080 ;
        RECT 31.380 16.500 31.640 16.760 ;
        RECT 31.380 16.180 31.640 16.440 ;
        RECT 32.960 19.380 33.220 19.640 ;
        RECT 32.960 19.060 33.220 19.320 ;
        RECT 32.960 18.740 33.220 19.000 ;
        RECT 32.960 18.420 33.220 18.680 ;
        RECT 32.960 18.100 33.220 18.360 ;
        RECT 32.960 17.780 33.220 18.040 ;
        RECT 32.960 17.460 33.220 17.720 ;
        RECT 32.960 17.140 33.220 17.400 ;
        RECT 32.960 16.820 33.220 17.080 ;
        RECT 32.960 16.500 33.220 16.760 ;
        RECT 32.960 16.180 33.220 16.440 ;
        RECT 34.540 19.380 34.800 19.640 ;
        RECT 34.540 19.060 34.800 19.320 ;
        RECT 34.540 18.740 34.800 19.000 ;
        RECT 34.540 18.420 34.800 18.680 ;
        RECT 34.540 18.100 34.800 18.360 ;
        RECT 34.540 17.780 34.800 18.040 ;
        RECT 34.540 17.460 34.800 17.720 ;
        RECT 34.540 17.140 34.800 17.400 ;
        RECT 34.540 16.820 34.800 17.080 ;
        RECT 34.540 16.500 34.800 16.760 ;
        RECT 34.540 16.180 34.800 16.440 ;
        RECT 36.120 19.380 36.380 19.640 ;
        RECT 36.120 19.060 36.380 19.320 ;
        RECT 36.120 18.740 36.380 19.000 ;
        RECT 36.120 18.420 36.380 18.680 ;
        RECT 36.120 18.100 36.380 18.360 ;
        RECT 36.120 17.780 36.380 18.040 ;
        RECT 36.120 17.460 36.380 17.720 ;
        RECT 36.120 17.140 36.380 17.400 ;
        RECT 36.120 16.820 36.380 17.080 ;
        RECT 36.120 16.500 36.380 16.760 ;
        RECT 36.120 16.180 36.380 16.440 ;
        RECT 37.700 19.380 37.960 19.640 ;
        RECT 37.700 19.060 37.960 19.320 ;
        RECT 37.700 18.740 37.960 19.000 ;
        RECT 37.700 18.420 37.960 18.680 ;
        RECT 37.700 18.100 37.960 18.360 ;
        RECT 37.700 17.780 37.960 18.040 ;
        RECT 37.700 17.460 37.960 17.720 ;
        RECT 37.700 17.140 37.960 17.400 ;
        RECT 37.700 16.820 37.960 17.080 ;
        RECT 37.700 16.500 37.960 16.760 ;
        RECT 37.700 16.180 37.960 16.440 ;
        RECT 39.280 19.380 39.540 19.640 ;
        RECT 39.280 19.060 39.540 19.320 ;
        RECT 39.280 18.740 39.540 19.000 ;
        RECT 39.280 18.420 39.540 18.680 ;
        RECT 39.280 18.100 39.540 18.360 ;
        RECT 39.280 17.780 39.540 18.040 ;
        RECT 39.280 17.460 39.540 17.720 ;
        RECT 39.280 17.140 39.540 17.400 ;
        RECT 39.280 16.820 39.540 17.080 ;
        RECT 39.280 16.500 39.540 16.760 ;
        RECT 39.280 16.180 39.540 16.440 ;
        RECT 40.860 19.380 41.120 19.640 ;
        RECT 40.860 19.060 41.120 19.320 ;
        RECT 40.860 18.740 41.120 19.000 ;
        RECT 40.860 18.420 41.120 18.680 ;
        RECT 40.860 18.100 41.120 18.360 ;
        RECT 40.860 17.780 41.120 18.040 ;
        RECT 40.860 17.460 41.120 17.720 ;
        RECT 40.860 17.140 41.120 17.400 ;
        RECT 40.860 16.820 41.120 17.080 ;
        RECT 40.860 16.500 41.120 16.760 ;
        RECT 40.860 16.180 41.120 16.440 ;
        RECT 42.440 19.380 42.700 19.640 ;
        RECT 42.440 19.060 42.700 19.320 ;
        RECT 42.440 18.740 42.700 19.000 ;
        RECT 42.440 18.420 42.700 18.680 ;
        RECT 42.440 18.100 42.700 18.360 ;
        RECT 42.440 17.780 42.700 18.040 ;
        RECT 42.440 17.460 42.700 17.720 ;
        RECT 42.440 17.140 42.700 17.400 ;
        RECT 42.440 16.820 42.700 17.080 ;
        RECT 42.440 16.500 42.700 16.760 ;
        RECT 42.440 16.180 42.700 16.440 ;
        RECT 44.020 19.380 44.280 19.640 ;
        RECT 44.020 19.060 44.280 19.320 ;
        RECT 44.020 18.740 44.280 19.000 ;
        RECT 44.020 18.420 44.280 18.680 ;
        RECT 44.020 18.100 44.280 18.360 ;
        RECT 44.020 17.780 44.280 18.040 ;
        RECT 44.020 17.460 44.280 17.720 ;
        RECT 44.020 17.140 44.280 17.400 ;
        RECT 44.020 16.820 44.280 17.080 ;
        RECT 44.020 16.500 44.280 16.760 ;
        RECT 44.020 16.180 44.280 16.440 ;
        RECT 45.600 19.380 45.860 19.640 ;
        RECT 45.600 19.060 45.860 19.320 ;
        RECT 45.600 18.740 45.860 19.000 ;
        RECT 45.600 18.420 45.860 18.680 ;
        RECT 45.600 18.100 45.860 18.360 ;
        RECT 45.600 17.780 45.860 18.040 ;
        RECT 45.600 17.460 45.860 17.720 ;
        RECT 45.600 17.140 45.860 17.400 ;
        RECT 45.600 16.820 45.860 17.080 ;
        RECT 45.600 16.500 45.860 16.760 ;
        RECT 45.600 16.180 45.860 16.440 ;
        RECT 47.180 19.380 47.440 19.640 ;
        RECT 47.180 19.060 47.440 19.320 ;
        RECT 47.180 18.740 47.440 19.000 ;
        RECT 47.180 18.420 47.440 18.680 ;
        RECT 47.180 18.100 47.440 18.360 ;
        RECT 47.180 17.780 47.440 18.040 ;
        RECT 47.180 17.460 47.440 17.720 ;
        RECT 47.180 17.140 47.440 17.400 ;
        RECT 47.180 16.820 47.440 17.080 ;
        RECT 47.180 16.500 47.440 16.760 ;
        RECT 47.180 16.180 47.440 16.440 ;
        RECT 51.100 16.335 52.000 19.475 ;
      LAYER met2 ;
        RECT -16.420 34.630 68.480 43.765 ;
        RECT 2.765 25.620 51.805 34.630 ;
        RECT 2.680 22.745 51.925 25.620 ;
        RECT 24.145 19.750 52.255 19.795 ;
        RECT 0.715 18.170 20.605 18.750 ;
        RECT 24.145 16.030 68.500 19.750 ;
        RECT -16.420 -35.805 68.480 -26.670 ;
      LAYER via2 ;
        RECT -15.885 35.185 -8.405 43.065 ;
        RECT 5.210 37.945 54.690 41.825 ;
        RECT 60.365 35.195 67.845 43.075 ;
        RECT 60.195 16.275 68.075 19.355 ;
        RECT -15.745 -35.075 -9.065 -27.595 ;
        RECT 60.640 -34.880 67.320 -27.400 ;
      LAYER met3 ;
        RECT -16.420 -35.805 -7.860 43.765 ;
        RECT 4.495 37.365 55.245 42.515 ;
        RECT 59.920 -35.805 68.480 43.765 ;
      LAYER via3 ;
        RECT 5.190 37.925 54.710 41.845 ;
      LAYER met4 ;
        RECT 4.495 35.755 55.245 42.515 ;
        RECT -4.375 27.260 57.910 35.755 ;
        RECT -4.375 26.145 25.235 27.260 ;
        RECT 28.300 26.145 57.910 27.260 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 141.518402 ;
    PORT
      LAYER pwell ;
        RECT 0.235 10.035 21.425 11.520 ;
        RECT 0.235 2.225 1.765 10.035 ;
        RECT 19.895 2.225 21.425 10.035 ;
        RECT 0.235 0.740 21.425 2.225 ;
        RECT 0.405 -0.985 14.300 0.145 ;
        RECT 0.405 -13.610 1.870 -0.985 ;
        RECT 12.835 -13.610 14.300 -0.985 ;
        RECT 0.405 -14.720 14.300 -13.610 ;
        RECT 0.405 -14.730 1.870 -14.720 ;
      LAYER li1 ;
        RECT 0.365 10.165 21.295 11.390 ;
        RECT 0.365 2.095 1.635 10.165 ;
        RECT 20.025 2.095 21.295 10.165 ;
        RECT 0.365 0.870 21.295 2.095 ;
        RECT 0.535 -0.855 19.655 0.870 ;
        RECT 0.535 -13.740 1.740 -0.855 ;
        RECT 4.020 -12.415 4.190 -1.875 ;
        RECT 5.600 -12.415 5.770 -1.875 ;
        RECT 7.180 -12.415 7.350 -1.875 ;
        RECT 8.760 -12.415 8.930 -1.875 ;
        RECT 10.340 -12.415 10.510 -1.875 ;
        RECT 12.270 -13.740 19.655 -0.855 ;
        RECT 0.535 -14.590 19.655 -13.740 ;
        RECT 0.535 -14.600 1.740 -14.590 ;
        RECT 12.270 -19.855 19.655 -14.590 ;
      LAYER mcon ;
        RECT 0.675 -6.785 1.565 -5.895 ;
        RECT 4.020 -2.190 4.190 -2.020 ;
        RECT 4.020 -2.550 4.190 -2.380 ;
        RECT 4.020 -2.910 4.190 -2.740 ;
        RECT 4.020 -3.270 4.190 -3.100 ;
        RECT 4.020 -3.630 4.190 -3.460 ;
        RECT 4.020 -3.990 4.190 -3.820 ;
        RECT 4.020 -4.350 4.190 -4.180 ;
        RECT 4.020 -4.710 4.190 -4.540 ;
        RECT 4.020 -5.070 4.190 -4.900 ;
        RECT 4.020 -5.430 4.190 -5.260 ;
        RECT 4.020 -5.790 4.190 -5.620 ;
        RECT 4.020 -6.150 4.190 -5.980 ;
        RECT 4.020 -6.510 4.190 -6.340 ;
        RECT 4.020 -6.870 4.190 -6.700 ;
        RECT 4.020 -7.230 4.190 -7.060 ;
        RECT 4.020 -7.590 4.190 -7.420 ;
        RECT 4.020 -7.950 4.190 -7.780 ;
        RECT 4.020 -8.310 4.190 -8.140 ;
        RECT 4.020 -8.670 4.190 -8.500 ;
        RECT 4.020 -9.030 4.190 -8.860 ;
        RECT 4.020 -9.390 4.190 -9.220 ;
        RECT 4.020 -9.750 4.190 -9.580 ;
        RECT 4.020 -10.110 4.190 -9.940 ;
        RECT 4.020 -10.470 4.190 -10.300 ;
        RECT 4.020 -10.830 4.190 -10.660 ;
        RECT 4.020 -11.190 4.190 -11.020 ;
        RECT 4.020 -11.550 4.190 -11.380 ;
        RECT 4.020 -11.910 4.190 -11.740 ;
        RECT 4.020 -12.270 4.190 -12.100 ;
        RECT 5.600 -2.190 5.770 -2.020 ;
        RECT 5.600 -2.550 5.770 -2.380 ;
        RECT 5.600 -2.910 5.770 -2.740 ;
        RECT 5.600 -3.270 5.770 -3.100 ;
        RECT 5.600 -3.630 5.770 -3.460 ;
        RECT 5.600 -3.990 5.770 -3.820 ;
        RECT 5.600 -4.350 5.770 -4.180 ;
        RECT 5.600 -4.710 5.770 -4.540 ;
        RECT 5.600 -5.070 5.770 -4.900 ;
        RECT 5.600 -5.430 5.770 -5.260 ;
        RECT 5.600 -5.790 5.770 -5.620 ;
        RECT 5.600 -6.150 5.770 -5.980 ;
        RECT 5.600 -6.510 5.770 -6.340 ;
        RECT 5.600 -6.870 5.770 -6.700 ;
        RECT 5.600 -7.230 5.770 -7.060 ;
        RECT 5.600 -7.590 5.770 -7.420 ;
        RECT 5.600 -7.950 5.770 -7.780 ;
        RECT 5.600 -8.310 5.770 -8.140 ;
        RECT 5.600 -8.670 5.770 -8.500 ;
        RECT 5.600 -9.030 5.770 -8.860 ;
        RECT 5.600 -9.390 5.770 -9.220 ;
        RECT 5.600 -9.750 5.770 -9.580 ;
        RECT 5.600 -10.110 5.770 -9.940 ;
        RECT 5.600 -10.470 5.770 -10.300 ;
        RECT 5.600 -10.830 5.770 -10.660 ;
        RECT 5.600 -11.190 5.770 -11.020 ;
        RECT 5.600 -11.550 5.770 -11.380 ;
        RECT 5.600 -11.910 5.770 -11.740 ;
        RECT 5.600 -12.270 5.770 -12.100 ;
        RECT 7.180 -2.190 7.350 -2.020 ;
        RECT 7.180 -2.550 7.350 -2.380 ;
        RECT 7.180 -2.910 7.350 -2.740 ;
        RECT 7.180 -3.270 7.350 -3.100 ;
        RECT 7.180 -3.630 7.350 -3.460 ;
        RECT 7.180 -3.990 7.350 -3.820 ;
        RECT 7.180 -4.350 7.350 -4.180 ;
        RECT 7.180 -4.710 7.350 -4.540 ;
        RECT 7.180 -5.070 7.350 -4.900 ;
        RECT 7.180 -5.430 7.350 -5.260 ;
        RECT 7.180 -5.790 7.350 -5.620 ;
        RECT 7.180 -6.150 7.350 -5.980 ;
        RECT 7.180 -6.510 7.350 -6.340 ;
        RECT 7.180 -6.870 7.350 -6.700 ;
        RECT 7.180 -7.230 7.350 -7.060 ;
        RECT 7.180 -7.590 7.350 -7.420 ;
        RECT 7.180 -7.950 7.350 -7.780 ;
        RECT 7.180 -8.310 7.350 -8.140 ;
        RECT 7.180 -8.670 7.350 -8.500 ;
        RECT 7.180 -9.030 7.350 -8.860 ;
        RECT 7.180 -9.390 7.350 -9.220 ;
        RECT 7.180 -9.750 7.350 -9.580 ;
        RECT 7.180 -10.110 7.350 -9.940 ;
        RECT 7.180 -10.470 7.350 -10.300 ;
        RECT 7.180 -10.830 7.350 -10.660 ;
        RECT 7.180 -11.190 7.350 -11.020 ;
        RECT 7.180 -11.550 7.350 -11.380 ;
        RECT 7.180 -11.910 7.350 -11.740 ;
        RECT 7.180 -12.270 7.350 -12.100 ;
        RECT 8.760 -2.190 8.930 -2.020 ;
        RECT 8.760 -2.550 8.930 -2.380 ;
        RECT 8.760 -2.910 8.930 -2.740 ;
        RECT 8.760 -3.270 8.930 -3.100 ;
        RECT 8.760 -3.630 8.930 -3.460 ;
        RECT 8.760 -3.990 8.930 -3.820 ;
        RECT 8.760 -4.350 8.930 -4.180 ;
        RECT 8.760 -4.710 8.930 -4.540 ;
        RECT 8.760 -5.070 8.930 -4.900 ;
        RECT 8.760 -5.430 8.930 -5.260 ;
        RECT 8.760 -5.790 8.930 -5.620 ;
        RECT 8.760 -6.150 8.930 -5.980 ;
        RECT 8.760 -6.510 8.930 -6.340 ;
        RECT 8.760 -6.870 8.930 -6.700 ;
        RECT 8.760 -7.230 8.930 -7.060 ;
        RECT 8.760 -7.590 8.930 -7.420 ;
        RECT 8.760 -7.950 8.930 -7.780 ;
        RECT 8.760 -8.310 8.930 -8.140 ;
        RECT 8.760 -8.670 8.930 -8.500 ;
        RECT 8.760 -9.030 8.930 -8.860 ;
        RECT 8.760 -9.390 8.930 -9.220 ;
        RECT 8.760 -9.750 8.930 -9.580 ;
        RECT 8.760 -10.110 8.930 -9.940 ;
        RECT 8.760 -10.470 8.930 -10.300 ;
        RECT 8.760 -10.830 8.930 -10.660 ;
        RECT 8.760 -11.190 8.930 -11.020 ;
        RECT 8.760 -11.550 8.930 -11.380 ;
        RECT 8.760 -11.910 8.930 -11.740 ;
        RECT 8.760 -12.270 8.930 -12.100 ;
        RECT 10.340 -2.190 10.510 -2.020 ;
        RECT 10.340 -2.550 10.510 -2.380 ;
        RECT 10.340 -2.910 10.510 -2.740 ;
        RECT 10.340 -3.270 10.510 -3.100 ;
        RECT 10.340 -3.630 10.510 -3.460 ;
        RECT 10.340 -3.990 10.510 -3.820 ;
        RECT 10.340 -4.350 10.510 -4.180 ;
        RECT 10.340 -4.710 10.510 -4.540 ;
        RECT 10.340 -5.070 10.510 -4.900 ;
        RECT 10.340 -5.430 10.510 -5.260 ;
        RECT 10.340 -5.790 10.510 -5.620 ;
        RECT 10.340 -6.150 10.510 -5.980 ;
        RECT 10.340 -6.510 10.510 -6.340 ;
        RECT 10.340 -6.870 10.510 -6.700 ;
        RECT 10.340 -7.230 10.510 -7.060 ;
        RECT 10.340 -7.590 10.510 -7.420 ;
        RECT 10.340 -7.950 10.510 -7.780 ;
        RECT 10.340 -8.310 10.510 -8.140 ;
        RECT 10.340 -8.670 10.510 -8.500 ;
        RECT 10.340 -9.030 10.510 -8.860 ;
        RECT 10.340 -9.390 10.510 -9.220 ;
        RECT 10.340 -9.750 10.510 -9.580 ;
        RECT 10.340 -10.110 10.510 -9.940 ;
        RECT 10.340 -10.470 10.510 -10.300 ;
        RECT 10.340 -10.830 10.510 -10.660 ;
        RECT 10.340 -11.190 10.510 -11.020 ;
        RECT 10.340 -11.550 10.510 -11.380 ;
        RECT 10.340 -11.910 10.510 -11.740 ;
        RECT 10.340 -12.270 10.510 -12.100 ;
        RECT 13.120 -6.790 14.010 -5.900 ;
        RECT 12.555 -19.550 19.205 -17.580 ;
      LAYER met1 ;
        RECT 3.990 -5.660 4.220 -1.895 ;
        RECT 5.570 -5.660 5.800 -1.895 ;
        RECT 7.150 -5.660 7.380 -1.895 ;
        RECT 8.730 -5.660 8.960 -1.895 ;
        RECT 10.310 -5.660 10.540 -1.895 ;
        RECT 0.535 -7.010 1.740 -5.660 ;
        RECT 3.945 -7.015 4.265 -5.660 ;
        RECT 5.525 -7.015 5.845 -5.660 ;
        RECT 7.105 -7.015 7.425 -5.660 ;
        RECT 8.685 -7.015 9.005 -5.660 ;
        RECT 10.265 -7.015 10.585 -5.660 ;
        RECT 12.965 -7.010 14.170 -5.660 ;
        RECT 3.990 -12.395 4.220 -7.015 ;
        RECT 5.570 -12.395 5.800 -7.015 ;
        RECT 7.150 -12.395 7.380 -7.015 ;
        RECT 8.730 -12.395 8.960 -7.015 ;
        RECT 10.310 -12.395 10.540 -7.015 ;
        RECT 12.270 -19.855 19.655 -17.165 ;
      LAYER via ;
        RECT 0.670 -6.790 1.570 -5.890 ;
        RECT 3.975 -5.990 4.235 -5.730 ;
        RECT 3.975 -6.310 4.235 -6.050 ;
        RECT 3.975 -6.630 4.235 -6.370 ;
        RECT 3.975 -6.950 4.235 -6.690 ;
        RECT 5.555 -5.990 5.815 -5.730 ;
        RECT 5.555 -6.310 5.815 -6.050 ;
        RECT 5.555 -6.630 5.815 -6.370 ;
        RECT 5.555 -6.950 5.815 -6.690 ;
        RECT 7.135 -5.990 7.395 -5.730 ;
        RECT 7.135 -6.310 7.395 -6.050 ;
        RECT 7.135 -6.630 7.395 -6.370 ;
        RECT 7.135 -6.950 7.395 -6.690 ;
        RECT 8.715 -5.990 8.975 -5.730 ;
        RECT 8.715 -6.310 8.975 -6.050 ;
        RECT 8.715 -6.630 8.975 -6.370 ;
        RECT 8.715 -6.950 8.975 -6.690 ;
        RECT 10.295 -5.990 10.555 -5.730 ;
        RECT 10.295 -6.310 10.555 -6.050 ;
        RECT 10.295 -6.630 10.555 -6.370 ;
        RECT 10.295 -6.950 10.555 -6.690 ;
        RECT 13.115 -6.795 14.015 -5.895 ;
        RECT 12.550 -19.655 19.210 -17.475 ;
      LAYER met2 ;
        RECT -31.050 45.320 84.480 57.360 ;
        RECT 0.535 -7.010 14.170 -5.660 ;
        RECT 12.270 -19.855 19.655 -17.165 ;
        RECT -31.050 -50.020 84.480 -37.980 ;
      LAYER via2 ;
        RECT -30.595 45.710 -20.715 56.790 ;
        RECT -7.845 46.100 -5.965 56.380 ;
        RECT 59.380 46.510 66.460 55.590 ;
        RECT 73.995 45.930 83.875 56.610 ;
        RECT 12.540 -19.705 19.220 -17.425 ;
        RECT -30.520 -49.310 -20.640 -39.030 ;
        RECT 12.950 -49.155 18.830 -38.875 ;
        RECT 74.310 -48.855 83.390 -38.975 ;
      LAYER met3 ;
        RECT -31.050 45.320 -20.040 57.370 ;
        RECT -8.500 45.320 -5.205 57.360 ;
        RECT 58.600 45.320 67.430 57.360 ;
        RECT -31.050 -50.020 -19.985 45.320 ;
        RECT -5.565 25.450 25.930 36.450 ;
        RECT 27.605 25.450 59.100 36.450 ;
        RECT 12.270 -50.020 19.655 -17.165 ;
        RECT 73.375 -50.020 84.480 57.360 ;
      LAYER via3 ;
        RECT -7.865 46.080 -5.945 56.400 ;
        RECT 59.560 46.490 66.280 55.610 ;
        RECT -5.465 35.990 -5.145 36.310 ;
        RECT -5.465 35.590 -5.145 35.910 ;
        RECT -5.465 35.190 -5.145 35.510 ;
        RECT -5.465 34.790 -5.145 35.110 ;
        RECT -5.465 34.390 -5.145 34.710 ;
        RECT -5.465 33.990 -5.145 34.310 ;
        RECT -5.465 33.590 -5.145 33.910 ;
        RECT -5.465 33.190 -5.145 33.510 ;
        RECT -5.465 32.790 -5.145 33.110 ;
        RECT -5.465 32.390 -5.145 32.710 ;
        RECT -5.465 31.990 -5.145 32.310 ;
        RECT -5.465 31.590 -5.145 31.910 ;
        RECT -5.465 31.190 -5.145 31.510 ;
        RECT -5.465 30.790 -5.145 31.110 ;
        RECT -5.465 30.390 -5.145 30.710 ;
        RECT -5.465 29.990 -5.145 30.310 ;
        RECT -5.465 29.590 -5.145 29.910 ;
        RECT -5.465 29.190 -5.145 29.510 ;
        RECT -5.465 28.790 -5.145 29.110 ;
        RECT -5.465 28.390 -5.145 28.710 ;
        RECT -5.465 27.990 -5.145 28.310 ;
        RECT -5.465 27.590 -5.145 27.910 ;
        RECT -5.465 27.190 -5.145 27.510 ;
        RECT -5.465 26.790 -5.145 27.110 ;
        RECT -5.465 26.390 -5.145 26.710 ;
        RECT -5.465 25.990 -5.145 26.310 ;
        RECT -5.465 25.590 -5.145 25.910 ;
        RECT 58.680 35.990 59.000 36.310 ;
        RECT 58.680 35.590 59.000 35.910 ;
        RECT 58.680 35.190 59.000 35.510 ;
        RECT 58.680 34.790 59.000 35.110 ;
        RECT 58.680 34.390 59.000 34.710 ;
        RECT 58.680 33.990 59.000 34.310 ;
        RECT 58.680 33.590 59.000 33.910 ;
        RECT 58.680 33.190 59.000 33.510 ;
        RECT 58.680 32.790 59.000 33.110 ;
        RECT 58.680 32.390 59.000 32.710 ;
        RECT 58.680 31.990 59.000 32.310 ;
        RECT 58.680 31.590 59.000 31.910 ;
        RECT 58.680 31.190 59.000 31.510 ;
        RECT 58.680 30.790 59.000 31.110 ;
        RECT 58.680 30.390 59.000 30.710 ;
        RECT 58.680 29.990 59.000 30.310 ;
        RECT 58.680 29.590 59.000 29.910 ;
        RECT 58.680 29.190 59.000 29.510 ;
        RECT 58.680 28.790 59.000 29.110 ;
        RECT 58.680 28.390 59.000 28.710 ;
        RECT 58.680 27.990 59.000 28.310 ;
        RECT 58.680 27.590 59.000 27.910 ;
        RECT 58.680 27.190 59.000 27.510 ;
        RECT 58.680 26.790 59.000 27.110 ;
        RECT 58.680 26.390 59.000 26.710 ;
        RECT 58.680 25.990 59.000 26.310 ;
        RECT 58.680 25.590 59.000 25.910 ;
      LAYER met4 ;
        RECT -8.500 36.390 -5.205 57.360 ;
        RECT -8.500 25.515 -5.065 36.390 ;
        RECT -5.545 25.510 -5.065 25.515 ;
        RECT 58.600 25.510 67.430 57.360 ;
    END
  END VSS
  PIN VO
    ANTENNADIFFAREA 65.713997 ;
    PORT
      LAYER li1 ;
        RECT 29.055 5.725 29.225 19.965 ;
        RECT 30.635 5.725 30.805 19.965 ;
        RECT 32.215 5.725 32.385 19.965 ;
        RECT 33.795 5.725 33.965 19.965 ;
        RECT 35.375 5.725 35.545 19.965 ;
        RECT 36.955 5.725 37.125 19.965 ;
        RECT 38.535 5.725 38.705 19.965 ;
        RECT 40.115 5.725 40.285 19.965 ;
        RECT 41.695 5.725 41.865 19.965 ;
        RECT 43.275 5.725 43.445 19.965 ;
        RECT 44.855 5.725 45.025 19.965 ;
        RECT 46.435 5.725 46.605 19.965 ;
        RECT 48.015 5.725 48.185 19.965 ;
        RECT 3.230 -12.415 3.400 -1.875 ;
        RECT 6.390 -12.415 6.560 -1.875 ;
        RECT 9.550 -12.415 9.720 -1.875 ;
        RECT 11.130 -12.415 11.300 -1.875 ;
      LAYER mcon ;
        RECT 29.055 19.600 29.225 19.770 ;
        RECT 29.055 19.240 29.225 19.410 ;
        RECT 29.055 18.880 29.225 19.050 ;
        RECT 29.055 18.520 29.225 18.690 ;
        RECT 29.055 18.160 29.225 18.330 ;
        RECT 29.055 17.800 29.225 17.970 ;
        RECT 29.055 17.440 29.225 17.610 ;
        RECT 29.055 17.080 29.225 17.250 ;
        RECT 29.055 16.720 29.225 16.890 ;
        RECT 29.055 16.360 29.225 16.530 ;
        RECT 29.055 16.000 29.225 16.170 ;
        RECT 29.055 15.640 29.225 15.810 ;
        RECT 29.055 15.280 29.225 15.450 ;
        RECT 29.055 14.920 29.225 15.090 ;
        RECT 29.055 14.560 29.225 14.730 ;
        RECT 29.055 14.200 29.225 14.370 ;
        RECT 29.055 13.840 29.225 14.010 ;
        RECT 29.055 13.480 29.225 13.650 ;
        RECT 29.055 13.120 29.225 13.290 ;
        RECT 29.055 12.760 29.225 12.930 ;
        RECT 29.055 12.400 29.225 12.570 ;
        RECT 29.055 12.040 29.225 12.210 ;
        RECT 29.055 11.680 29.225 11.850 ;
        RECT 29.055 11.320 29.225 11.490 ;
        RECT 29.055 10.960 29.225 11.130 ;
        RECT 29.055 10.600 29.225 10.770 ;
        RECT 29.055 10.240 29.225 10.410 ;
        RECT 29.055 9.880 29.225 10.050 ;
        RECT 29.055 9.520 29.225 9.690 ;
        RECT 29.055 9.160 29.225 9.330 ;
        RECT 29.055 8.800 29.225 8.970 ;
        RECT 29.055 8.440 29.225 8.610 ;
        RECT 29.055 8.080 29.225 8.250 ;
        RECT 29.055 7.720 29.225 7.890 ;
        RECT 29.055 7.360 29.225 7.530 ;
        RECT 29.055 7.000 29.225 7.170 ;
        RECT 29.055 6.640 29.225 6.810 ;
        RECT 29.055 6.280 29.225 6.450 ;
        RECT 29.055 5.920 29.225 6.090 ;
        RECT 30.635 19.600 30.805 19.770 ;
        RECT 30.635 19.240 30.805 19.410 ;
        RECT 30.635 18.880 30.805 19.050 ;
        RECT 30.635 18.520 30.805 18.690 ;
        RECT 30.635 18.160 30.805 18.330 ;
        RECT 30.635 17.800 30.805 17.970 ;
        RECT 30.635 17.440 30.805 17.610 ;
        RECT 30.635 17.080 30.805 17.250 ;
        RECT 30.635 16.720 30.805 16.890 ;
        RECT 30.635 16.360 30.805 16.530 ;
        RECT 30.635 16.000 30.805 16.170 ;
        RECT 30.635 15.640 30.805 15.810 ;
        RECT 30.635 15.280 30.805 15.450 ;
        RECT 30.635 14.920 30.805 15.090 ;
        RECT 30.635 14.560 30.805 14.730 ;
        RECT 30.635 14.200 30.805 14.370 ;
        RECT 30.635 13.840 30.805 14.010 ;
        RECT 30.635 13.480 30.805 13.650 ;
        RECT 30.635 13.120 30.805 13.290 ;
        RECT 30.635 12.760 30.805 12.930 ;
        RECT 30.635 12.400 30.805 12.570 ;
        RECT 30.635 12.040 30.805 12.210 ;
        RECT 30.635 11.680 30.805 11.850 ;
        RECT 30.635 11.320 30.805 11.490 ;
        RECT 30.635 10.960 30.805 11.130 ;
        RECT 30.635 10.600 30.805 10.770 ;
        RECT 30.635 10.240 30.805 10.410 ;
        RECT 30.635 9.880 30.805 10.050 ;
        RECT 30.635 9.520 30.805 9.690 ;
        RECT 30.635 9.160 30.805 9.330 ;
        RECT 30.635 8.800 30.805 8.970 ;
        RECT 30.635 8.440 30.805 8.610 ;
        RECT 30.635 8.080 30.805 8.250 ;
        RECT 30.635 7.720 30.805 7.890 ;
        RECT 30.635 7.360 30.805 7.530 ;
        RECT 30.635 7.000 30.805 7.170 ;
        RECT 30.635 6.640 30.805 6.810 ;
        RECT 30.635 6.280 30.805 6.450 ;
        RECT 30.635 5.920 30.805 6.090 ;
        RECT 32.215 19.600 32.385 19.770 ;
        RECT 32.215 19.240 32.385 19.410 ;
        RECT 32.215 18.880 32.385 19.050 ;
        RECT 32.215 18.520 32.385 18.690 ;
        RECT 32.215 18.160 32.385 18.330 ;
        RECT 32.215 17.800 32.385 17.970 ;
        RECT 32.215 17.440 32.385 17.610 ;
        RECT 32.215 17.080 32.385 17.250 ;
        RECT 32.215 16.720 32.385 16.890 ;
        RECT 32.215 16.360 32.385 16.530 ;
        RECT 32.215 16.000 32.385 16.170 ;
        RECT 32.215 15.640 32.385 15.810 ;
        RECT 32.215 15.280 32.385 15.450 ;
        RECT 32.215 14.920 32.385 15.090 ;
        RECT 32.215 14.560 32.385 14.730 ;
        RECT 32.215 14.200 32.385 14.370 ;
        RECT 32.215 13.840 32.385 14.010 ;
        RECT 32.215 13.480 32.385 13.650 ;
        RECT 32.215 13.120 32.385 13.290 ;
        RECT 32.215 12.760 32.385 12.930 ;
        RECT 32.215 12.400 32.385 12.570 ;
        RECT 32.215 12.040 32.385 12.210 ;
        RECT 32.215 11.680 32.385 11.850 ;
        RECT 32.215 11.320 32.385 11.490 ;
        RECT 32.215 10.960 32.385 11.130 ;
        RECT 32.215 10.600 32.385 10.770 ;
        RECT 32.215 10.240 32.385 10.410 ;
        RECT 32.215 9.880 32.385 10.050 ;
        RECT 32.215 9.520 32.385 9.690 ;
        RECT 32.215 9.160 32.385 9.330 ;
        RECT 32.215 8.800 32.385 8.970 ;
        RECT 32.215 8.440 32.385 8.610 ;
        RECT 32.215 8.080 32.385 8.250 ;
        RECT 32.215 7.720 32.385 7.890 ;
        RECT 32.215 7.360 32.385 7.530 ;
        RECT 32.215 7.000 32.385 7.170 ;
        RECT 32.215 6.640 32.385 6.810 ;
        RECT 32.215 6.280 32.385 6.450 ;
        RECT 32.215 5.920 32.385 6.090 ;
        RECT 33.795 19.600 33.965 19.770 ;
        RECT 33.795 19.240 33.965 19.410 ;
        RECT 33.795 18.880 33.965 19.050 ;
        RECT 33.795 18.520 33.965 18.690 ;
        RECT 33.795 18.160 33.965 18.330 ;
        RECT 33.795 17.800 33.965 17.970 ;
        RECT 33.795 17.440 33.965 17.610 ;
        RECT 33.795 17.080 33.965 17.250 ;
        RECT 33.795 16.720 33.965 16.890 ;
        RECT 33.795 16.360 33.965 16.530 ;
        RECT 33.795 16.000 33.965 16.170 ;
        RECT 33.795 15.640 33.965 15.810 ;
        RECT 33.795 15.280 33.965 15.450 ;
        RECT 33.795 14.920 33.965 15.090 ;
        RECT 33.795 14.560 33.965 14.730 ;
        RECT 33.795 14.200 33.965 14.370 ;
        RECT 33.795 13.840 33.965 14.010 ;
        RECT 33.795 13.480 33.965 13.650 ;
        RECT 33.795 13.120 33.965 13.290 ;
        RECT 33.795 12.760 33.965 12.930 ;
        RECT 33.795 12.400 33.965 12.570 ;
        RECT 33.795 12.040 33.965 12.210 ;
        RECT 33.795 11.680 33.965 11.850 ;
        RECT 33.795 11.320 33.965 11.490 ;
        RECT 33.795 10.960 33.965 11.130 ;
        RECT 33.795 10.600 33.965 10.770 ;
        RECT 33.795 10.240 33.965 10.410 ;
        RECT 33.795 9.880 33.965 10.050 ;
        RECT 33.795 9.520 33.965 9.690 ;
        RECT 33.795 9.160 33.965 9.330 ;
        RECT 33.795 8.800 33.965 8.970 ;
        RECT 33.795 8.440 33.965 8.610 ;
        RECT 33.795 8.080 33.965 8.250 ;
        RECT 33.795 7.720 33.965 7.890 ;
        RECT 33.795 7.360 33.965 7.530 ;
        RECT 33.795 7.000 33.965 7.170 ;
        RECT 33.795 6.640 33.965 6.810 ;
        RECT 33.795 6.280 33.965 6.450 ;
        RECT 33.795 5.920 33.965 6.090 ;
        RECT 35.375 19.600 35.545 19.770 ;
        RECT 35.375 19.240 35.545 19.410 ;
        RECT 35.375 18.880 35.545 19.050 ;
        RECT 35.375 18.520 35.545 18.690 ;
        RECT 35.375 18.160 35.545 18.330 ;
        RECT 35.375 17.800 35.545 17.970 ;
        RECT 35.375 17.440 35.545 17.610 ;
        RECT 35.375 17.080 35.545 17.250 ;
        RECT 35.375 16.720 35.545 16.890 ;
        RECT 35.375 16.360 35.545 16.530 ;
        RECT 35.375 16.000 35.545 16.170 ;
        RECT 35.375 15.640 35.545 15.810 ;
        RECT 35.375 15.280 35.545 15.450 ;
        RECT 35.375 14.920 35.545 15.090 ;
        RECT 35.375 14.560 35.545 14.730 ;
        RECT 35.375 14.200 35.545 14.370 ;
        RECT 35.375 13.840 35.545 14.010 ;
        RECT 35.375 13.480 35.545 13.650 ;
        RECT 35.375 13.120 35.545 13.290 ;
        RECT 35.375 12.760 35.545 12.930 ;
        RECT 35.375 12.400 35.545 12.570 ;
        RECT 35.375 12.040 35.545 12.210 ;
        RECT 35.375 11.680 35.545 11.850 ;
        RECT 35.375 11.320 35.545 11.490 ;
        RECT 35.375 10.960 35.545 11.130 ;
        RECT 35.375 10.600 35.545 10.770 ;
        RECT 35.375 10.240 35.545 10.410 ;
        RECT 35.375 9.880 35.545 10.050 ;
        RECT 35.375 9.520 35.545 9.690 ;
        RECT 35.375 9.160 35.545 9.330 ;
        RECT 35.375 8.800 35.545 8.970 ;
        RECT 35.375 8.440 35.545 8.610 ;
        RECT 35.375 8.080 35.545 8.250 ;
        RECT 35.375 7.720 35.545 7.890 ;
        RECT 35.375 7.360 35.545 7.530 ;
        RECT 35.375 7.000 35.545 7.170 ;
        RECT 35.375 6.640 35.545 6.810 ;
        RECT 35.375 6.280 35.545 6.450 ;
        RECT 35.375 5.920 35.545 6.090 ;
        RECT 36.955 19.600 37.125 19.770 ;
        RECT 36.955 19.240 37.125 19.410 ;
        RECT 36.955 18.880 37.125 19.050 ;
        RECT 36.955 18.520 37.125 18.690 ;
        RECT 36.955 18.160 37.125 18.330 ;
        RECT 36.955 17.800 37.125 17.970 ;
        RECT 36.955 17.440 37.125 17.610 ;
        RECT 36.955 17.080 37.125 17.250 ;
        RECT 36.955 16.720 37.125 16.890 ;
        RECT 36.955 16.360 37.125 16.530 ;
        RECT 36.955 16.000 37.125 16.170 ;
        RECT 36.955 15.640 37.125 15.810 ;
        RECT 36.955 15.280 37.125 15.450 ;
        RECT 36.955 14.920 37.125 15.090 ;
        RECT 36.955 14.560 37.125 14.730 ;
        RECT 36.955 14.200 37.125 14.370 ;
        RECT 36.955 13.840 37.125 14.010 ;
        RECT 36.955 13.480 37.125 13.650 ;
        RECT 36.955 13.120 37.125 13.290 ;
        RECT 36.955 12.760 37.125 12.930 ;
        RECT 36.955 12.400 37.125 12.570 ;
        RECT 36.955 12.040 37.125 12.210 ;
        RECT 36.955 11.680 37.125 11.850 ;
        RECT 36.955 11.320 37.125 11.490 ;
        RECT 36.955 10.960 37.125 11.130 ;
        RECT 36.955 10.600 37.125 10.770 ;
        RECT 36.955 10.240 37.125 10.410 ;
        RECT 36.955 9.880 37.125 10.050 ;
        RECT 36.955 9.520 37.125 9.690 ;
        RECT 36.955 9.160 37.125 9.330 ;
        RECT 36.955 8.800 37.125 8.970 ;
        RECT 36.955 8.440 37.125 8.610 ;
        RECT 36.955 8.080 37.125 8.250 ;
        RECT 36.955 7.720 37.125 7.890 ;
        RECT 36.955 7.360 37.125 7.530 ;
        RECT 36.955 7.000 37.125 7.170 ;
        RECT 36.955 6.640 37.125 6.810 ;
        RECT 36.955 6.280 37.125 6.450 ;
        RECT 36.955 5.920 37.125 6.090 ;
        RECT 38.535 19.600 38.705 19.770 ;
        RECT 38.535 19.240 38.705 19.410 ;
        RECT 38.535 18.880 38.705 19.050 ;
        RECT 38.535 18.520 38.705 18.690 ;
        RECT 38.535 18.160 38.705 18.330 ;
        RECT 38.535 17.800 38.705 17.970 ;
        RECT 38.535 17.440 38.705 17.610 ;
        RECT 38.535 17.080 38.705 17.250 ;
        RECT 38.535 16.720 38.705 16.890 ;
        RECT 38.535 16.360 38.705 16.530 ;
        RECT 38.535 16.000 38.705 16.170 ;
        RECT 38.535 15.640 38.705 15.810 ;
        RECT 38.535 15.280 38.705 15.450 ;
        RECT 38.535 14.920 38.705 15.090 ;
        RECT 38.535 14.560 38.705 14.730 ;
        RECT 38.535 14.200 38.705 14.370 ;
        RECT 38.535 13.840 38.705 14.010 ;
        RECT 38.535 13.480 38.705 13.650 ;
        RECT 38.535 13.120 38.705 13.290 ;
        RECT 38.535 12.760 38.705 12.930 ;
        RECT 38.535 12.400 38.705 12.570 ;
        RECT 38.535 12.040 38.705 12.210 ;
        RECT 38.535 11.680 38.705 11.850 ;
        RECT 38.535 11.320 38.705 11.490 ;
        RECT 38.535 10.960 38.705 11.130 ;
        RECT 38.535 10.600 38.705 10.770 ;
        RECT 38.535 10.240 38.705 10.410 ;
        RECT 38.535 9.880 38.705 10.050 ;
        RECT 38.535 9.520 38.705 9.690 ;
        RECT 38.535 9.160 38.705 9.330 ;
        RECT 38.535 8.800 38.705 8.970 ;
        RECT 38.535 8.440 38.705 8.610 ;
        RECT 38.535 8.080 38.705 8.250 ;
        RECT 38.535 7.720 38.705 7.890 ;
        RECT 38.535 7.360 38.705 7.530 ;
        RECT 38.535 7.000 38.705 7.170 ;
        RECT 38.535 6.640 38.705 6.810 ;
        RECT 38.535 6.280 38.705 6.450 ;
        RECT 38.535 5.920 38.705 6.090 ;
        RECT 40.115 19.600 40.285 19.770 ;
        RECT 40.115 19.240 40.285 19.410 ;
        RECT 40.115 18.880 40.285 19.050 ;
        RECT 40.115 18.520 40.285 18.690 ;
        RECT 40.115 18.160 40.285 18.330 ;
        RECT 40.115 17.800 40.285 17.970 ;
        RECT 40.115 17.440 40.285 17.610 ;
        RECT 40.115 17.080 40.285 17.250 ;
        RECT 40.115 16.720 40.285 16.890 ;
        RECT 40.115 16.360 40.285 16.530 ;
        RECT 40.115 16.000 40.285 16.170 ;
        RECT 40.115 15.640 40.285 15.810 ;
        RECT 40.115 15.280 40.285 15.450 ;
        RECT 40.115 14.920 40.285 15.090 ;
        RECT 40.115 14.560 40.285 14.730 ;
        RECT 40.115 14.200 40.285 14.370 ;
        RECT 40.115 13.840 40.285 14.010 ;
        RECT 40.115 13.480 40.285 13.650 ;
        RECT 40.115 13.120 40.285 13.290 ;
        RECT 40.115 12.760 40.285 12.930 ;
        RECT 40.115 12.400 40.285 12.570 ;
        RECT 40.115 12.040 40.285 12.210 ;
        RECT 40.115 11.680 40.285 11.850 ;
        RECT 40.115 11.320 40.285 11.490 ;
        RECT 40.115 10.960 40.285 11.130 ;
        RECT 40.115 10.600 40.285 10.770 ;
        RECT 40.115 10.240 40.285 10.410 ;
        RECT 40.115 9.880 40.285 10.050 ;
        RECT 40.115 9.520 40.285 9.690 ;
        RECT 40.115 9.160 40.285 9.330 ;
        RECT 40.115 8.800 40.285 8.970 ;
        RECT 40.115 8.440 40.285 8.610 ;
        RECT 40.115 8.080 40.285 8.250 ;
        RECT 40.115 7.720 40.285 7.890 ;
        RECT 40.115 7.360 40.285 7.530 ;
        RECT 40.115 7.000 40.285 7.170 ;
        RECT 40.115 6.640 40.285 6.810 ;
        RECT 40.115 6.280 40.285 6.450 ;
        RECT 40.115 5.920 40.285 6.090 ;
        RECT 41.695 19.600 41.865 19.770 ;
        RECT 41.695 19.240 41.865 19.410 ;
        RECT 41.695 18.880 41.865 19.050 ;
        RECT 41.695 18.520 41.865 18.690 ;
        RECT 41.695 18.160 41.865 18.330 ;
        RECT 41.695 17.800 41.865 17.970 ;
        RECT 41.695 17.440 41.865 17.610 ;
        RECT 41.695 17.080 41.865 17.250 ;
        RECT 41.695 16.720 41.865 16.890 ;
        RECT 41.695 16.360 41.865 16.530 ;
        RECT 41.695 16.000 41.865 16.170 ;
        RECT 41.695 15.640 41.865 15.810 ;
        RECT 41.695 15.280 41.865 15.450 ;
        RECT 41.695 14.920 41.865 15.090 ;
        RECT 41.695 14.560 41.865 14.730 ;
        RECT 41.695 14.200 41.865 14.370 ;
        RECT 41.695 13.840 41.865 14.010 ;
        RECT 41.695 13.480 41.865 13.650 ;
        RECT 41.695 13.120 41.865 13.290 ;
        RECT 41.695 12.760 41.865 12.930 ;
        RECT 41.695 12.400 41.865 12.570 ;
        RECT 41.695 12.040 41.865 12.210 ;
        RECT 41.695 11.680 41.865 11.850 ;
        RECT 41.695 11.320 41.865 11.490 ;
        RECT 41.695 10.960 41.865 11.130 ;
        RECT 41.695 10.600 41.865 10.770 ;
        RECT 41.695 10.240 41.865 10.410 ;
        RECT 41.695 9.880 41.865 10.050 ;
        RECT 41.695 9.520 41.865 9.690 ;
        RECT 41.695 9.160 41.865 9.330 ;
        RECT 41.695 8.800 41.865 8.970 ;
        RECT 41.695 8.440 41.865 8.610 ;
        RECT 41.695 8.080 41.865 8.250 ;
        RECT 41.695 7.720 41.865 7.890 ;
        RECT 41.695 7.360 41.865 7.530 ;
        RECT 41.695 7.000 41.865 7.170 ;
        RECT 41.695 6.640 41.865 6.810 ;
        RECT 41.695 6.280 41.865 6.450 ;
        RECT 41.695 5.920 41.865 6.090 ;
        RECT 43.275 19.600 43.445 19.770 ;
        RECT 43.275 19.240 43.445 19.410 ;
        RECT 43.275 18.880 43.445 19.050 ;
        RECT 43.275 18.520 43.445 18.690 ;
        RECT 43.275 18.160 43.445 18.330 ;
        RECT 43.275 17.800 43.445 17.970 ;
        RECT 43.275 17.440 43.445 17.610 ;
        RECT 43.275 17.080 43.445 17.250 ;
        RECT 43.275 16.720 43.445 16.890 ;
        RECT 43.275 16.360 43.445 16.530 ;
        RECT 43.275 16.000 43.445 16.170 ;
        RECT 43.275 15.640 43.445 15.810 ;
        RECT 43.275 15.280 43.445 15.450 ;
        RECT 43.275 14.920 43.445 15.090 ;
        RECT 43.275 14.560 43.445 14.730 ;
        RECT 43.275 14.200 43.445 14.370 ;
        RECT 43.275 13.840 43.445 14.010 ;
        RECT 43.275 13.480 43.445 13.650 ;
        RECT 43.275 13.120 43.445 13.290 ;
        RECT 43.275 12.760 43.445 12.930 ;
        RECT 43.275 12.400 43.445 12.570 ;
        RECT 43.275 12.040 43.445 12.210 ;
        RECT 43.275 11.680 43.445 11.850 ;
        RECT 43.275 11.320 43.445 11.490 ;
        RECT 43.275 10.960 43.445 11.130 ;
        RECT 43.275 10.600 43.445 10.770 ;
        RECT 43.275 10.240 43.445 10.410 ;
        RECT 43.275 9.880 43.445 10.050 ;
        RECT 43.275 9.520 43.445 9.690 ;
        RECT 43.275 9.160 43.445 9.330 ;
        RECT 43.275 8.800 43.445 8.970 ;
        RECT 43.275 8.440 43.445 8.610 ;
        RECT 43.275 8.080 43.445 8.250 ;
        RECT 43.275 7.720 43.445 7.890 ;
        RECT 43.275 7.360 43.445 7.530 ;
        RECT 43.275 7.000 43.445 7.170 ;
        RECT 43.275 6.640 43.445 6.810 ;
        RECT 43.275 6.280 43.445 6.450 ;
        RECT 43.275 5.920 43.445 6.090 ;
        RECT 44.855 19.600 45.025 19.770 ;
        RECT 44.855 19.240 45.025 19.410 ;
        RECT 44.855 18.880 45.025 19.050 ;
        RECT 44.855 18.520 45.025 18.690 ;
        RECT 44.855 18.160 45.025 18.330 ;
        RECT 44.855 17.800 45.025 17.970 ;
        RECT 44.855 17.440 45.025 17.610 ;
        RECT 44.855 17.080 45.025 17.250 ;
        RECT 44.855 16.720 45.025 16.890 ;
        RECT 44.855 16.360 45.025 16.530 ;
        RECT 44.855 16.000 45.025 16.170 ;
        RECT 44.855 15.640 45.025 15.810 ;
        RECT 44.855 15.280 45.025 15.450 ;
        RECT 44.855 14.920 45.025 15.090 ;
        RECT 44.855 14.560 45.025 14.730 ;
        RECT 44.855 14.200 45.025 14.370 ;
        RECT 44.855 13.840 45.025 14.010 ;
        RECT 44.855 13.480 45.025 13.650 ;
        RECT 44.855 13.120 45.025 13.290 ;
        RECT 44.855 12.760 45.025 12.930 ;
        RECT 44.855 12.400 45.025 12.570 ;
        RECT 44.855 12.040 45.025 12.210 ;
        RECT 44.855 11.680 45.025 11.850 ;
        RECT 44.855 11.320 45.025 11.490 ;
        RECT 44.855 10.960 45.025 11.130 ;
        RECT 44.855 10.600 45.025 10.770 ;
        RECT 44.855 10.240 45.025 10.410 ;
        RECT 44.855 9.880 45.025 10.050 ;
        RECT 44.855 9.520 45.025 9.690 ;
        RECT 44.855 9.160 45.025 9.330 ;
        RECT 44.855 8.800 45.025 8.970 ;
        RECT 44.855 8.440 45.025 8.610 ;
        RECT 44.855 8.080 45.025 8.250 ;
        RECT 44.855 7.720 45.025 7.890 ;
        RECT 44.855 7.360 45.025 7.530 ;
        RECT 44.855 7.000 45.025 7.170 ;
        RECT 44.855 6.640 45.025 6.810 ;
        RECT 44.855 6.280 45.025 6.450 ;
        RECT 44.855 5.920 45.025 6.090 ;
        RECT 46.435 19.600 46.605 19.770 ;
        RECT 46.435 19.240 46.605 19.410 ;
        RECT 46.435 18.880 46.605 19.050 ;
        RECT 46.435 18.520 46.605 18.690 ;
        RECT 46.435 18.160 46.605 18.330 ;
        RECT 46.435 17.800 46.605 17.970 ;
        RECT 46.435 17.440 46.605 17.610 ;
        RECT 46.435 17.080 46.605 17.250 ;
        RECT 46.435 16.720 46.605 16.890 ;
        RECT 46.435 16.360 46.605 16.530 ;
        RECT 46.435 16.000 46.605 16.170 ;
        RECT 46.435 15.640 46.605 15.810 ;
        RECT 46.435 15.280 46.605 15.450 ;
        RECT 46.435 14.920 46.605 15.090 ;
        RECT 46.435 14.560 46.605 14.730 ;
        RECT 46.435 14.200 46.605 14.370 ;
        RECT 46.435 13.840 46.605 14.010 ;
        RECT 46.435 13.480 46.605 13.650 ;
        RECT 46.435 13.120 46.605 13.290 ;
        RECT 46.435 12.760 46.605 12.930 ;
        RECT 46.435 12.400 46.605 12.570 ;
        RECT 46.435 12.040 46.605 12.210 ;
        RECT 46.435 11.680 46.605 11.850 ;
        RECT 46.435 11.320 46.605 11.490 ;
        RECT 46.435 10.960 46.605 11.130 ;
        RECT 46.435 10.600 46.605 10.770 ;
        RECT 46.435 10.240 46.605 10.410 ;
        RECT 46.435 9.880 46.605 10.050 ;
        RECT 46.435 9.520 46.605 9.690 ;
        RECT 46.435 9.160 46.605 9.330 ;
        RECT 46.435 8.800 46.605 8.970 ;
        RECT 46.435 8.440 46.605 8.610 ;
        RECT 46.435 8.080 46.605 8.250 ;
        RECT 46.435 7.720 46.605 7.890 ;
        RECT 46.435 7.360 46.605 7.530 ;
        RECT 46.435 7.000 46.605 7.170 ;
        RECT 46.435 6.640 46.605 6.810 ;
        RECT 46.435 6.280 46.605 6.450 ;
        RECT 46.435 5.920 46.605 6.090 ;
        RECT 48.015 19.600 48.185 19.770 ;
        RECT 48.015 19.240 48.185 19.410 ;
        RECT 48.015 18.880 48.185 19.050 ;
        RECT 48.015 18.520 48.185 18.690 ;
        RECT 48.015 18.160 48.185 18.330 ;
        RECT 48.015 17.800 48.185 17.970 ;
        RECT 48.015 17.440 48.185 17.610 ;
        RECT 48.015 17.080 48.185 17.250 ;
        RECT 48.015 16.720 48.185 16.890 ;
        RECT 48.015 16.360 48.185 16.530 ;
        RECT 48.015 16.000 48.185 16.170 ;
        RECT 48.015 15.640 48.185 15.810 ;
        RECT 48.015 15.280 48.185 15.450 ;
        RECT 48.015 14.920 48.185 15.090 ;
        RECT 48.015 14.560 48.185 14.730 ;
        RECT 48.015 14.200 48.185 14.370 ;
        RECT 48.015 13.840 48.185 14.010 ;
        RECT 48.015 13.480 48.185 13.650 ;
        RECT 48.015 13.120 48.185 13.290 ;
        RECT 48.015 12.760 48.185 12.930 ;
        RECT 48.015 12.400 48.185 12.570 ;
        RECT 48.015 12.040 48.185 12.210 ;
        RECT 48.015 11.680 48.185 11.850 ;
        RECT 48.015 11.320 48.185 11.490 ;
        RECT 48.015 10.960 48.185 11.130 ;
        RECT 48.015 10.600 48.185 10.770 ;
        RECT 48.015 10.240 48.185 10.410 ;
        RECT 48.015 9.880 48.185 10.050 ;
        RECT 48.015 9.520 48.185 9.690 ;
        RECT 48.015 9.160 48.185 9.330 ;
        RECT 48.015 8.800 48.185 8.970 ;
        RECT 48.015 8.440 48.185 8.610 ;
        RECT 48.015 8.080 48.185 8.250 ;
        RECT 48.015 7.720 48.185 7.890 ;
        RECT 48.015 7.360 48.185 7.530 ;
        RECT 48.015 7.000 48.185 7.170 ;
        RECT 48.015 6.640 48.185 6.810 ;
        RECT 48.015 6.280 48.185 6.450 ;
        RECT 48.015 5.920 48.185 6.090 ;
        RECT 3.230 -2.190 3.400 -2.020 ;
        RECT 3.230 -2.550 3.400 -2.380 ;
        RECT 3.230 -2.910 3.400 -2.740 ;
        RECT 3.230 -3.270 3.400 -3.100 ;
        RECT 3.230 -3.630 3.400 -3.460 ;
        RECT 3.230 -3.990 3.400 -3.820 ;
        RECT 3.230 -4.350 3.400 -4.180 ;
        RECT 3.230 -4.710 3.400 -4.540 ;
        RECT 3.230 -5.070 3.400 -4.900 ;
        RECT 3.230 -5.430 3.400 -5.260 ;
        RECT 3.230 -5.790 3.400 -5.620 ;
        RECT 3.230 -6.150 3.400 -5.980 ;
        RECT 3.230 -6.510 3.400 -6.340 ;
        RECT 3.230 -6.870 3.400 -6.700 ;
        RECT 3.230 -7.230 3.400 -7.060 ;
        RECT 3.230 -7.590 3.400 -7.420 ;
        RECT 3.230 -7.950 3.400 -7.780 ;
        RECT 3.230 -8.310 3.400 -8.140 ;
        RECT 3.230 -8.670 3.400 -8.500 ;
        RECT 3.230 -9.030 3.400 -8.860 ;
        RECT 3.230 -9.390 3.400 -9.220 ;
        RECT 3.230 -9.750 3.400 -9.580 ;
        RECT 3.230 -10.110 3.400 -9.940 ;
        RECT 3.230 -10.470 3.400 -10.300 ;
        RECT 3.230 -10.830 3.400 -10.660 ;
        RECT 3.230 -11.190 3.400 -11.020 ;
        RECT 3.230 -11.550 3.400 -11.380 ;
        RECT 3.230 -11.910 3.400 -11.740 ;
        RECT 3.230 -12.270 3.400 -12.100 ;
        RECT 6.390 -2.190 6.560 -2.020 ;
        RECT 6.390 -2.550 6.560 -2.380 ;
        RECT 6.390 -2.910 6.560 -2.740 ;
        RECT 6.390 -3.270 6.560 -3.100 ;
        RECT 6.390 -3.630 6.560 -3.460 ;
        RECT 6.390 -3.990 6.560 -3.820 ;
        RECT 6.390 -4.350 6.560 -4.180 ;
        RECT 6.390 -4.710 6.560 -4.540 ;
        RECT 6.390 -5.070 6.560 -4.900 ;
        RECT 6.390 -5.430 6.560 -5.260 ;
        RECT 6.390 -5.790 6.560 -5.620 ;
        RECT 6.390 -6.150 6.560 -5.980 ;
        RECT 6.390 -6.510 6.560 -6.340 ;
        RECT 6.390 -6.870 6.560 -6.700 ;
        RECT 6.390 -7.230 6.560 -7.060 ;
        RECT 6.390 -7.590 6.560 -7.420 ;
        RECT 6.390 -7.950 6.560 -7.780 ;
        RECT 6.390 -8.310 6.560 -8.140 ;
        RECT 6.390 -8.670 6.560 -8.500 ;
        RECT 6.390 -9.030 6.560 -8.860 ;
        RECT 6.390 -9.390 6.560 -9.220 ;
        RECT 6.390 -9.750 6.560 -9.580 ;
        RECT 6.390 -10.110 6.560 -9.940 ;
        RECT 6.390 -10.470 6.560 -10.300 ;
        RECT 6.390 -10.830 6.560 -10.660 ;
        RECT 6.390 -11.190 6.560 -11.020 ;
        RECT 6.390 -11.550 6.560 -11.380 ;
        RECT 6.390 -11.910 6.560 -11.740 ;
        RECT 6.390 -12.270 6.560 -12.100 ;
        RECT 9.550 -2.190 9.720 -2.020 ;
        RECT 9.550 -2.550 9.720 -2.380 ;
        RECT 9.550 -2.910 9.720 -2.740 ;
        RECT 9.550 -3.270 9.720 -3.100 ;
        RECT 9.550 -3.630 9.720 -3.460 ;
        RECT 9.550 -3.990 9.720 -3.820 ;
        RECT 9.550 -4.350 9.720 -4.180 ;
        RECT 9.550 -4.710 9.720 -4.540 ;
        RECT 9.550 -5.070 9.720 -4.900 ;
        RECT 9.550 -5.430 9.720 -5.260 ;
        RECT 9.550 -5.790 9.720 -5.620 ;
        RECT 9.550 -6.150 9.720 -5.980 ;
        RECT 9.550 -6.510 9.720 -6.340 ;
        RECT 9.550 -6.870 9.720 -6.700 ;
        RECT 9.550 -7.230 9.720 -7.060 ;
        RECT 9.550 -7.590 9.720 -7.420 ;
        RECT 9.550 -7.950 9.720 -7.780 ;
        RECT 9.550 -8.310 9.720 -8.140 ;
        RECT 9.550 -8.670 9.720 -8.500 ;
        RECT 9.550 -9.030 9.720 -8.860 ;
        RECT 9.550 -9.390 9.720 -9.220 ;
        RECT 9.550 -9.750 9.720 -9.580 ;
        RECT 9.550 -10.110 9.720 -9.940 ;
        RECT 9.550 -10.470 9.720 -10.300 ;
        RECT 9.550 -10.830 9.720 -10.660 ;
        RECT 9.550 -11.190 9.720 -11.020 ;
        RECT 9.550 -11.550 9.720 -11.380 ;
        RECT 9.550 -11.910 9.720 -11.740 ;
        RECT 9.550 -12.270 9.720 -12.100 ;
        RECT 11.130 -2.190 11.300 -2.020 ;
        RECT 11.130 -2.550 11.300 -2.380 ;
        RECT 11.130 -2.910 11.300 -2.740 ;
        RECT 11.130 -3.270 11.300 -3.100 ;
        RECT 11.130 -3.630 11.300 -3.460 ;
        RECT 11.130 -3.990 11.300 -3.820 ;
        RECT 11.130 -4.350 11.300 -4.180 ;
        RECT 11.130 -4.710 11.300 -4.540 ;
        RECT 11.130 -5.070 11.300 -4.900 ;
        RECT 11.130 -5.430 11.300 -5.260 ;
        RECT 11.130 -5.790 11.300 -5.620 ;
        RECT 11.130 -6.150 11.300 -5.980 ;
        RECT 11.130 -6.510 11.300 -6.340 ;
        RECT 11.130 -6.870 11.300 -6.700 ;
        RECT 11.130 -7.230 11.300 -7.060 ;
        RECT 11.130 -7.590 11.300 -7.420 ;
        RECT 11.130 -7.950 11.300 -7.780 ;
        RECT 11.130 -8.310 11.300 -8.140 ;
        RECT 11.130 -8.670 11.300 -8.500 ;
        RECT 11.130 -9.030 11.300 -8.860 ;
        RECT 11.130 -9.390 11.300 -9.220 ;
        RECT 11.130 -9.750 11.300 -9.580 ;
        RECT 11.130 -10.110 11.300 -9.940 ;
        RECT 11.130 -10.470 11.300 -10.300 ;
        RECT 11.130 -10.830 11.300 -10.660 ;
        RECT 11.130 -11.190 11.300 -11.020 ;
        RECT 11.130 -11.550 11.300 -11.380 ;
        RECT 11.130 -11.910 11.300 -11.740 ;
        RECT 11.130 -12.270 11.300 -12.100 ;
      LAYER met1 ;
        RECT 29.025 10.615 29.255 19.945 ;
        RECT 30.605 10.615 30.835 19.945 ;
        RECT 32.185 10.615 32.415 19.945 ;
        RECT 33.765 10.615 33.995 19.945 ;
        RECT 35.345 10.615 35.575 19.945 ;
        RECT 36.925 10.615 37.155 19.945 ;
        RECT 38.505 10.615 38.735 19.945 ;
        RECT 40.085 10.615 40.315 19.945 ;
        RECT 41.665 10.615 41.895 19.945 ;
        RECT 43.245 10.615 43.475 19.945 ;
        RECT 44.825 10.615 45.055 19.945 ;
        RECT 46.405 10.615 46.635 19.945 ;
        RECT 47.985 10.615 48.215 19.945 ;
        RECT 28.980 6.860 29.300 10.615 ;
        RECT 30.560 6.860 30.880 10.615 ;
        RECT 32.140 6.860 32.460 10.615 ;
        RECT 33.720 6.860 34.040 10.615 ;
        RECT 35.300 6.860 35.620 10.615 ;
        RECT 36.880 6.860 37.200 10.615 ;
        RECT 38.460 6.860 38.780 10.615 ;
        RECT 40.040 6.860 40.360 10.615 ;
        RECT 41.620 6.860 41.940 10.615 ;
        RECT 43.200 6.860 43.520 10.615 ;
        RECT 44.780 6.860 45.100 10.615 ;
        RECT 46.360 6.860 46.680 10.615 ;
        RECT 47.940 6.860 48.260 10.615 ;
        RECT 29.025 5.745 29.255 6.860 ;
        RECT 30.605 5.745 30.835 6.860 ;
        RECT 32.185 5.745 32.415 6.860 ;
        RECT 33.765 5.745 33.995 6.860 ;
        RECT 35.345 5.745 35.575 6.860 ;
        RECT 36.925 5.745 37.155 6.860 ;
        RECT 38.505 5.745 38.735 6.860 ;
        RECT 40.085 5.745 40.315 6.860 ;
        RECT 41.665 5.745 41.895 6.860 ;
        RECT 43.245 5.745 43.475 6.860 ;
        RECT 44.825 5.745 45.055 6.860 ;
        RECT 46.405 5.745 46.635 6.860 ;
        RECT 47.985 5.745 48.215 6.860 ;
        RECT 3.200 -11.115 3.430 -1.895 ;
        RECT 6.360 -11.115 6.590 -1.895 ;
        RECT 9.520 -11.115 9.750 -1.895 ;
        RECT 11.100 -11.115 11.330 -1.895 ;
        RECT 3.155 -11.950 3.475 -11.115 ;
        RECT 6.315 -11.950 6.635 -11.115 ;
        RECT 9.475 -11.950 9.795 -11.115 ;
        RECT 11.055 -11.950 11.375 -11.115 ;
        RECT 3.200 -12.395 3.430 -11.950 ;
        RECT 6.360 -12.395 6.590 -11.950 ;
        RECT 9.520 -12.395 9.750 -11.950 ;
        RECT 11.100 -12.395 11.330 -11.950 ;
      LAYER via ;
        RECT 29.010 10.185 29.270 10.445 ;
        RECT 29.010 9.865 29.270 10.125 ;
        RECT 29.010 9.545 29.270 9.805 ;
        RECT 29.010 9.225 29.270 9.485 ;
        RECT 29.010 8.905 29.270 9.165 ;
        RECT 29.010 8.585 29.270 8.845 ;
        RECT 29.010 8.265 29.270 8.525 ;
        RECT 29.010 7.945 29.270 8.205 ;
        RECT 29.010 7.625 29.270 7.885 ;
        RECT 29.010 7.305 29.270 7.565 ;
        RECT 29.010 6.985 29.270 7.245 ;
        RECT 30.590 10.185 30.850 10.445 ;
        RECT 30.590 9.865 30.850 10.125 ;
        RECT 30.590 9.545 30.850 9.805 ;
        RECT 30.590 9.225 30.850 9.485 ;
        RECT 30.590 8.905 30.850 9.165 ;
        RECT 30.590 8.585 30.850 8.845 ;
        RECT 30.590 8.265 30.850 8.525 ;
        RECT 30.590 7.945 30.850 8.205 ;
        RECT 30.590 7.625 30.850 7.885 ;
        RECT 30.590 7.305 30.850 7.565 ;
        RECT 30.590 6.985 30.850 7.245 ;
        RECT 32.170 10.185 32.430 10.445 ;
        RECT 32.170 9.865 32.430 10.125 ;
        RECT 32.170 9.545 32.430 9.805 ;
        RECT 32.170 9.225 32.430 9.485 ;
        RECT 32.170 8.905 32.430 9.165 ;
        RECT 32.170 8.585 32.430 8.845 ;
        RECT 32.170 8.265 32.430 8.525 ;
        RECT 32.170 7.945 32.430 8.205 ;
        RECT 32.170 7.625 32.430 7.885 ;
        RECT 32.170 7.305 32.430 7.565 ;
        RECT 32.170 6.985 32.430 7.245 ;
        RECT 33.750 10.185 34.010 10.445 ;
        RECT 33.750 9.865 34.010 10.125 ;
        RECT 33.750 9.545 34.010 9.805 ;
        RECT 33.750 9.225 34.010 9.485 ;
        RECT 33.750 8.905 34.010 9.165 ;
        RECT 33.750 8.585 34.010 8.845 ;
        RECT 33.750 8.265 34.010 8.525 ;
        RECT 33.750 7.945 34.010 8.205 ;
        RECT 33.750 7.625 34.010 7.885 ;
        RECT 33.750 7.305 34.010 7.565 ;
        RECT 33.750 6.985 34.010 7.245 ;
        RECT 35.330 10.185 35.590 10.445 ;
        RECT 35.330 9.865 35.590 10.125 ;
        RECT 35.330 9.545 35.590 9.805 ;
        RECT 35.330 9.225 35.590 9.485 ;
        RECT 35.330 8.905 35.590 9.165 ;
        RECT 35.330 8.585 35.590 8.845 ;
        RECT 35.330 8.265 35.590 8.525 ;
        RECT 35.330 7.945 35.590 8.205 ;
        RECT 35.330 7.625 35.590 7.885 ;
        RECT 35.330 7.305 35.590 7.565 ;
        RECT 35.330 6.985 35.590 7.245 ;
        RECT 36.910 10.185 37.170 10.445 ;
        RECT 36.910 9.865 37.170 10.125 ;
        RECT 36.910 9.545 37.170 9.805 ;
        RECT 36.910 9.225 37.170 9.485 ;
        RECT 36.910 8.905 37.170 9.165 ;
        RECT 36.910 8.585 37.170 8.845 ;
        RECT 36.910 8.265 37.170 8.525 ;
        RECT 36.910 7.945 37.170 8.205 ;
        RECT 36.910 7.625 37.170 7.885 ;
        RECT 36.910 7.305 37.170 7.565 ;
        RECT 36.910 6.985 37.170 7.245 ;
        RECT 38.490 10.185 38.750 10.445 ;
        RECT 38.490 9.865 38.750 10.125 ;
        RECT 38.490 9.545 38.750 9.805 ;
        RECT 38.490 9.225 38.750 9.485 ;
        RECT 38.490 8.905 38.750 9.165 ;
        RECT 38.490 8.585 38.750 8.845 ;
        RECT 38.490 8.265 38.750 8.525 ;
        RECT 38.490 7.945 38.750 8.205 ;
        RECT 38.490 7.625 38.750 7.885 ;
        RECT 38.490 7.305 38.750 7.565 ;
        RECT 38.490 6.985 38.750 7.245 ;
        RECT 40.070 10.185 40.330 10.445 ;
        RECT 40.070 9.865 40.330 10.125 ;
        RECT 40.070 9.545 40.330 9.805 ;
        RECT 40.070 9.225 40.330 9.485 ;
        RECT 40.070 8.905 40.330 9.165 ;
        RECT 40.070 8.585 40.330 8.845 ;
        RECT 40.070 8.265 40.330 8.525 ;
        RECT 40.070 7.945 40.330 8.205 ;
        RECT 40.070 7.625 40.330 7.885 ;
        RECT 40.070 7.305 40.330 7.565 ;
        RECT 40.070 6.985 40.330 7.245 ;
        RECT 41.650 10.185 41.910 10.445 ;
        RECT 41.650 9.865 41.910 10.125 ;
        RECT 41.650 9.545 41.910 9.805 ;
        RECT 41.650 9.225 41.910 9.485 ;
        RECT 41.650 8.905 41.910 9.165 ;
        RECT 41.650 8.585 41.910 8.845 ;
        RECT 41.650 8.265 41.910 8.525 ;
        RECT 41.650 7.945 41.910 8.205 ;
        RECT 41.650 7.625 41.910 7.885 ;
        RECT 41.650 7.305 41.910 7.565 ;
        RECT 41.650 6.985 41.910 7.245 ;
        RECT 43.230 10.185 43.490 10.445 ;
        RECT 43.230 9.865 43.490 10.125 ;
        RECT 43.230 9.545 43.490 9.805 ;
        RECT 43.230 9.225 43.490 9.485 ;
        RECT 43.230 8.905 43.490 9.165 ;
        RECT 43.230 8.585 43.490 8.845 ;
        RECT 43.230 8.265 43.490 8.525 ;
        RECT 43.230 7.945 43.490 8.205 ;
        RECT 43.230 7.625 43.490 7.885 ;
        RECT 43.230 7.305 43.490 7.565 ;
        RECT 43.230 6.985 43.490 7.245 ;
        RECT 44.810 10.185 45.070 10.445 ;
        RECT 44.810 9.865 45.070 10.125 ;
        RECT 44.810 9.545 45.070 9.805 ;
        RECT 44.810 9.225 45.070 9.485 ;
        RECT 44.810 8.905 45.070 9.165 ;
        RECT 44.810 8.585 45.070 8.845 ;
        RECT 44.810 8.265 45.070 8.525 ;
        RECT 44.810 7.945 45.070 8.205 ;
        RECT 44.810 7.625 45.070 7.885 ;
        RECT 44.810 7.305 45.070 7.565 ;
        RECT 44.810 6.985 45.070 7.245 ;
        RECT 46.390 10.185 46.650 10.445 ;
        RECT 46.390 9.865 46.650 10.125 ;
        RECT 46.390 9.545 46.650 9.805 ;
        RECT 46.390 9.225 46.650 9.485 ;
        RECT 46.390 8.905 46.650 9.165 ;
        RECT 46.390 8.585 46.650 8.845 ;
        RECT 46.390 8.265 46.650 8.525 ;
        RECT 46.390 7.945 46.650 8.205 ;
        RECT 46.390 7.625 46.650 7.885 ;
        RECT 46.390 7.305 46.650 7.565 ;
        RECT 46.390 6.985 46.650 7.245 ;
        RECT 47.970 10.185 48.230 10.445 ;
        RECT 47.970 9.865 48.230 10.125 ;
        RECT 47.970 9.545 48.230 9.805 ;
        RECT 47.970 9.225 48.230 9.485 ;
        RECT 47.970 8.905 48.230 9.165 ;
        RECT 47.970 8.585 48.230 8.845 ;
        RECT 47.970 8.265 48.230 8.525 ;
        RECT 47.970 7.945 48.230 8.205 ;
        RECT 47.970 7.625 48.230 7.885 ;
        RECT 47.970 7.305 48.230 7.565 ;
        RECT 47.970 6.985 48.230 7.245 ;
        RECT 3.185 -11.505 3.445 -11.245 ;
        RECT 3.185 -11.825 3.445 -11.565 ;
        RECT 6.345 -11.505 6.605 -11.245 ;
        RECT 6.345 -11.825 6.605 -11.565 ;
        RECT 9.505 -11.505 9.765 -11.245 ;
        RECT 9.505 -11.825 9.765 -11.565 ;
        RECT 11.085 -11.505 11.345 -11.245 ;
        RECT 11.085 -11.825 11.345 -11.565 ;
      LAYER met2 ;
        RECT 28.205 10.595 48.245 10.615 ;
        RECT 28.205 6.860 55.115 10.595 ;
        RECT 10.540 -11.115 59.325 -8.180 ;
        RECT 3.155 -11.945 59.325 -11.115 ;
      LAYER via2 ;
        RECT 53.335 7.160 54.815 10.240 ;
        RECT 53.525 -11.365 58.605 -8.685 ;
      LAYER met3 ;
        RECT 53.120 6.860 55.115 10.595 ;
        RECT 27.625 -8.180 53.120 0.365 ;
        RECT 27.625 -11.945 59.325 -8.180 ;
        RECT 27.625 -24.635 53.120 -11.945 ;
      LAYER via3 ;
        RECT 53.515 7.140 54.635 10.260 ;
        RECT 52.700 -0.095 53.020 0.225 ;
        RECT 52.700 -0.495 53.020 -0.175 ;
        RECT 52.700 -0.895 53.020 -0.575 ;
        RECT 52.700 -1.295 53.020 -0.975 ;
        RECT 52.700 -1.695 53.020 -1.375 ;
        RECT 52.700 -2.095 53.020 -1.775 ;
        RECT 52.700 -2.495 53.020 -2.175 ;
        RECT 52.700 -2.895 53.020 -2.575 ;
        RECT 52.700 -3.295 53.020 -2.975 ;
        RECT 52.700 -3.695 53.020 -3.375 ;
        RECT 52.700 -4.095 53.020 -3.775 ;
        RECT 52.700 -4.495 53.020 -4.175 ;
        RECT 52.700 -4.895 53.020 -4.575 ;
        RECT 52.700 -5.295 53.020 -4.975 ;
        RECT 52.700 -5.695 53.020 -5.375 ;
        RECT 52.700 -6.095 53.020 -5.775 ;
        RECT 52.700 -6.495 53.020 -6.175 ;
        RECT 52.700 -6.895 53.020 -6.575 ;
        RECT 52.700 -7.295 53.020 -6.975 ;
        RECT 52.700 -7.695 53.020 -7.375 ;
        RECT 52.700 -8.095 53.020 -7.775 ;
        RECT 52.700 -8.495 53.020 -8.175 ;
        RECT 52.700 -8.895 53.020 -8.575 ;
        RECT 52.700 -9.295 53.020 -8.975 ;
        RECT 52.700 -9.695 53.020 -9.375 ;
        RECT 52.700 -10.095 53.020 -9.775 ;
        RECT 52.700 -10.495 53.020 -10.175 ;
        RECT 52.700 -10.895 53.020 -10.575 ;
        RECT 52.700 -11.295 53.020 -10.975 ;
        RECT 52.700 -11.695 53.020 -11.375 ;
        RECT 53.705 -11.385 58.425 -8.665 ;
        RECT 52.700 -12.095 53.020 -11.775 ;
        RECT 52.700 -12.495 53.020 -12.175 ;
        RECT 52.700 -12.895 53.020 -12.575 ;
        RECT 52.700 -13.295 53.020 -12.975 ;
        RECT 52.700 -13.695 53.020 -13.375 ;
        RECT 52.700 -14.095 53.020 -13.775 ;
        RECT 52.700 -14.495 53.020 -14.175 ;
        RECT 52.700 -14.895 53.020 -14.575 ;
        RECT 52.700 -15.295 53.020 -14.975 ;
        RECT 52.700 -15.695 53.020 -15.375 ;
        RECT 52.700 -16.095 53.020 -15.775 ;
        RECT 52.700 -16.495 53.020 -16.175 ;
        RECT 52.700 -16.895 53.020 -16.575 ;
        RECT 52.700 -17.295 53.020 -16.975 ;
        RECT 52.700 -17.695 53.020 -17.375 ;
        RECT 52.700 -18.095 53.020 -17.775 ;
        RECT 52.700 -18.495 53.020 -18.175 ;
        RECT 52.700 -18.895 53.020 -18.575 ;
        RECT 52.700 -19.295 53.020 -18.975 ;
        RECT 52.700 -19.695 53.020 -19.375 ;
        RECT 52.700 -20.095 53.020 -19.775 ;
        RECT 52.700 -20.495 53.020 -20.175 ;
        RECT 52.700 -20.895 53.020 -20.575 ;
        RECT 52.700 -21.295 53.020 -20.975 ;
        RECT 52.700 -21.695 53.020 -21.375 ;
        RECT 52.700 -22.095 53.020 -21.775 ;
        RECT 52.700 -22.495 53.020 -22.175 ;
        RECT 52.700 -22.895 53.020 -22.575 ;
        RECT 52.700 -23.295 53.020 -22.975 ;
        RECT 52.700 -23.695 53.020 -23.375 ;
        RECT 52.700 -24.095 53.020 -23.775 ;
        RECT 52.700 -24.495 53.020 -24.175 ;
      LAYER met4 ;
        RECT 53.120 4.975 60.155 10.605 ;
        RECT 53.120 0.305 105.020 4.975 ;
        RECT 52.620 -4.600 105.020 0.305 ;
        RECT 52.620 -8.180 55.115 -4.600 ;
        RECT 58.060 -7.120 105.020 -4.600 ;
        RECT 52.620 -11.945 59.325 -8.180 ;
        RECT 52.620 -24.575 55.115 -11.945 ;
    END
  END VO
  OBS
      LAYER pwell ;
        RECT 2.180 3.505 18.530 8.765 ;
        RECT 3.040 -12.525 11.490 -1.765 ;
      LAYER li1 ;
        RECT 2.920 21.910 18.430 22.230 ;
        RECT 2.690 15.550 2.860 21.590 ;
        RECT 4.270 15.550 4.440 21.590 ;
        RECT 5.850 15.550 6.020 21.590 ;
        RECT 7.430 15.550 7.600 21.590 ;
        RECT 9.010 15.550 9.180 21.590 ;
        RECT 10.590 15.550 10.760 21.590 ;
        RECT 12.170 15.550 12.340 21.590 ;
        RECT 13.750 15.550 13.920 21.590 ;
        RECT 15.330 15.550 15.500 21.590 ;
        RECT 16.910 15.550 17.080 21.590 ;
        RECT 18.490 15.550 18.660 21.590 ;
        RECT 28.495 20.285 47.955 20.605 ;
        RECT 2.920 14.910 18.430 15.230 ;
        RECT 2.370 3.615 2.540 8.655 ;
        RECT 3.160 3.615 3.330 8.655 ;
        RECT 3.950 3.615 4.120 8.655 ;
        RECT 4.740 3.615 4.910 8.655 ;
        RECT 5.530 3.615 5.700 8.655 ;
        RECT 6.320 3.615 6.490 8.655 ;
        RECT 7.110 3.615 7.280 8.655 ;
        RECT 7.900 3.615 8.070 8.655 ;
        RECT 8.690 3.615 8.860 8.655 ;
        RECT 9.480 3.615 9.650 8.655 ;
        RECT 10.270 3.615 10.440 8.655 ;
        RECT 11.060 3.615 11.230 8.655 ;
        RECT 11.850 3.615 12.020 8.655 ;
        RECT 12.640 3.615 12.810 8.655 ;
        RECT 13.430 3.615 13.600 8.655 ;
        RECT 14.220 3.615 14.390 8.655 ;
        RECT 15.010 3.615 15.180 8.655 ;
        RECT 15.800 3.615 15.970 8.655 ;
        RECT 16.590 3.615 16.760 8.655 ;
        RECT 17.380 3.615 17.550 8.655 ;
        RECT 18.170 3.615 18.340 8.655 ;
        RECT 28.495 5.085 47.955 5.405 ;
        RECT 4.810 -12.415 4.980 -1.875 ;
      LAYER mcon ;
        RECT 3.165 21.990 3.335 22.160 ;
        RECT 3.525 21.990 3.695 22.160 ;
        RECT 3.885 21.990 4.055 22.160 ;
        RECT 4.245 21.990 4.415 22.160 ;
        RECT 4.605 21.990 4.775 22.160 ;
        RECT 4.965 21.990 5.135 22.160 ;
        RECT 5.325 21.990 5.495 22.160 ;
        RECT 5.685 21.990 5.855 22.160 ;
        RECT 6.045 21.990 6.215 22.160 ;
        RECT 6.405 21.990 6.575 22.160 ;
        RECT 6.765 21.990 6.935 22.160 ;
        RECT 7.125 21.990 7.295 22.160 ;
        RECT 7.485 21.990 7.655 22.160 ;
        RECT 7.845 21.990 8.015 22.160 ;
        RECT 8.205 21.990 8.375 22.160 ;
        RECT 8.565 21.990 8.735 22.160 ;
        RECT 8.925 21.990 9.095 22.160 ;
        RECT 9.285 21.990 9.455 22.160 ;
        RECT 9.645 21.990 9.815 22.160 ;
        RECT 10.005 21.990 10.175 22.160 ;
        RECT 10.365 21.990 10.535 22.160 ;
        RECT 10.725 21.990 10.895 22.160 ;
        RECT 11.085 21.990 11.255 22.160 ;
        RECT 11.445 21.990 11.615 22.160 ;
        RECT 11.805 21.990 11.975 22.160 ;
        RECT 12.165 21.990 12.335 22.160 ;
        RECT 12.525 21.990 12.695 22.160 ;
        RECT 12.885 21.990 13.055 22.160 ;
        RECT 13.245 21.990 13.415 22.160 ;
        RECT 13.605 21.990 13.775 22.160 ;
        RECT 13.965 21.990 14.135 22.160 ;
        RECT 14.325 21.990 14.495 22.160 ;
        RECT 14.685 21.990 14.855 22.160 ;
        RECT 15.045 21.990 15.215 22.160 ;
        RECT 15.405 21.990 15.575 22.160 ;
        RECT 15.765 21.990 15.935 22.160 ;
        RECT 16.125 21.990 16.295 22.160 ;
        RECT 16.485 21.990 16.655 22.160 ;
        RECT 16.845 21.990 17.015 22.160 ;
        RECT 17.205 21.990 17.375 22.160 ;
        RECT 17.565 21.990 17.735 22.160 ;
        RECT 17.925 21.990 18.095 22.160 ;
        RECT 2.690 21.185 2.860 21.355 ;
        RECT 2.690 20.825 2.860 20.995 ;
        RECT 2.690 20.465 2.860 20.635 ;
        RECT 2.690 20.105 2.860 20.275 ;
        RECT 2.690 19.745 2.860 19.915 ;
        RECT 2.690 19.385 2.860 19.555 ;
        RECT 2.690 19.025 2.860 19.195 ;
        RECT 2.690 18.665 2.860 18.835 ;
        RECT 2.690 18.305 2.860 18.475 ;
        RECT 2.690 17.945 2.860 18.115 ;
        RECT 2.690 17.585 2.860 17.755 ;
        RECT 2.690 17.225 2.860 17.395 ;
        RECT 2.690 16.865 2.860 17.035 ;
        RECT 2.690 16.505 2.860 16.675 ;
        RECT 2.690 16.145 2.860 16.315 ;
        RECT 2.690 15.785 2.860 15.955 ;
        RECT 4.270 21.185 4.440 21.355 ;
        RECT 4.270 20.825 4.440 20.995 ;
        RECT 4.270 20.465 4.440 20.635 ;
        RECT 4.270 20.105 4.440 20.275 ;
        RECT 4.270 19.745 4.440 19.915 ;
        RECT 4.270 19.385 4.440 19.555 ;
        RECT 4.270 19.025 4.440 19.195 ;
        RECT 4.270 18.665 4.440 18.835 ;
        RECT 4.270 18.305 4.440 18.475 ;
        RECT 4.270 17.945 4.440 18.115 ;
        RECT 4.270 17.585 4.440 17.755 ;
        RECT 4.270 17.225 4.440 17.395 ;
        RECT 4.270 16.865 4.440 17.035 ;
        RECT 4.270 16.505 4.440 16.675 ;
        RECT 4.270 16.145 4.440 16.315 ;
        RECT 4.270 15.785 4.440 15.955 ;
        RECT 5.850 21.185 6.020 21.355 ;
        RECT 5.850 20.825 6.020 20.995 ;
        RECT 5.850 20.465 6.020 20.635 ;
        RECT 5.850 20.105 6.020 20.275 ;
        RECT 5.850 19.745 6.020 19.915 ;
        RECT 5.850 19.385 6.020 19.555 ;
        RECT 5.850 19.025 6.020 19.195 ;
        RECT 5.850 18.665 6.020 18.835 ;
        RECT 5.850 18.305 6.020 18.475 ;
        RECT 5.850 17.945 6.020 18.115 ;
        RECT 5.850 17.585 6.020 17.755 ;
        RECT 5.850 17.225 6.020 17.395 ;
        RECT 5.850 16.865 6.020 17.035 ;
        RECT 5.850 16.505 6.020 16.675 ;
        RECT 5.850 16.145 6.020 16.315 ;
        RECT 5.850 15.785 6.020 15.955 ;
        RECT 7.430 21.185 7.600 21.355 ;
        RECT 7.430 20.825 7.600 20.995 ;
        RECT 7.430 20.465 7.600 20.635 ;
        RECT 7.430 20.105 7.600 20.275 ;
        RECT 7.430 19.745 7.600 19.915 ;
        RECT 7.430 19.385 7.600 19.555 ;
        RECT 7.430 19.025 7.600 19.195 ;
        RECT 7.430 18.665 7.600 18.835 ;
        RECT 7.430 18.305 7.600 18.475 ;
        RECT 7.430 17.945 7.600 18.115 ;
        RECT 7.430 17.585 7.600 17.755 ;
        RECT 7.430 17.225 7.600 17.395 ;
        RECT 7.430 16.865 7.600 17.035 ;
        RECT 7.430 16.505 7.600 16.675 ;
        RECT 7.430 16.145 7.600 16.315 ;
        RECT 7.430 15.785 7.600 15.955 ;
        RECT 9.010 21.185 9.180 21.355 ;
        RECT 9.010 20.825 9.180 20.995 ;
        RECT 9.010 20.465 9.180 20.635 ;
        RECT 9.010 20.105 9.180 20.275 ;
        RECT 9.010 19.745 9.180 19.915 ;
        RECT 9.010 19.385 9.180 19.555 ;
        RECT 9.010 19.025 9.180 19.195 ;
        RECT 9.010 18.665 9.180 18.835 ;
        RECT 9.010 18.305 9.180 18.475 ;
        RECT 9.010 17.945 9.180 18.115 ;
        RECT 9.010 17.585 9.180 17.755 ;
        RECT 9.010 17.225 9.180 17.395 ;
        RECT 9.010 16.865 9.180 17.035 ;
        RECT 9.010 16.505 9.180 16.675 ;
        RECT 9.010 16.145 9.180 16.315 ;
        RECT 9.010 15.785 9.180 15.955 ;
        RECT 10.590 21.185 10.760 21.355 ;
        RECT 10.590 20.825 10.760 20.995 ;
        RECT 10.590 20.465 10.760 20.635 ;
        RECT 10.590 20.105 10.760 20.275 ;
        RECT 10.590 19.745 10.760 19.915 ;
        RECT 10.590 19.385 10.760 19.555 ;
        RECT 10.590 19.025 10.760 19.195 ;
        RECT 10.590 18.665 10.760 18.835 ;
        RECT 10.590 18.305 10.760 18.475 ;
        RECT 10.590 17.945 10.760 18.115 ;
        RECT 10.590 17.585 10.760 17.755 ;
        RECT 10.590 17.225 10.760 17.395 ;
        RECT 10.590 16.865 10.760 17.035 ;
        RECT 10.590 16.505 10.760 16.675 ;
        RECT 10.590 16.145 10.760 16.315 ;
        RECT 10.590 15.785 10.760 15.955 ;
        RECT 12.170 21.185 12.340 21.355 ;
        RECT 12.170 20.825 12.340 20.995 ;
        RECT 12.170 20.465 12.340 20.635 ;
        RECT 12.170 20.105 12.340 20.275 ;
        RECT 12.170 19.745 12.340 19.915 ;
        RECT 12.170 19.385 12.340 19.555 ;
        RECT 12.170 19.025 12.340 19.195 ;
        RECT 12.170 18.665 12.340 18.835 ;
        RECT 12.170 18.305 12.340 18.475 ;
        RECT 12.170 17.945 12.340 18.115 ;
        RECT 12.170 17.585 12.340 17.755 ;
        RECT 12.170 17.225 12.340 17.395 ;
        RECT 12.170 16.865 12.340 17.035 ;
        RECT 12.170 16.505 12.340 16.675 ;
        RECT 12.170 16.145 12.340 16.315 ;
        RECT 12.170 15.785 12.340 15.955 ;
        RECT 13.750 21.185 13.920 21.355 ;
        RECT 13.750 20.825 13.920 20.995 ;
        RECT 13.750 20.465 13.920 20.635 ;
        RECT 13.750 20.105 13.920 20.275 ;
        RECT 13.750 19.745 13.920 19.915 ;
        RECT 13.750 19.385 13.920 19.555 ;
        RECT 13.750 19.025 13.920 19.195 ;
        RECT 13.750 18.665 13.920 18.835 ;
        RECT 13.750 18.305 13.920 18.475 ;
        RECT 13.750 17.945 13.920 18.115 ;
        RECT 13.750 17.585 13.920 17.755 ;
        RECT 13.750 17.225 13.920 17.395 ;
        RECT 13.750 16.865 13.920 17.035 ;
        RECT 13.750 16.505 13.920 16.675 ;
        RECT 13.750 16.145 13.920 16.315 ;
        RECT 13.750 15.785 13.920 15.955 ;
        RECT 15.330 21.185 15.500 21.355 ;
        RECT 15.330 20.825 15.500 20.995 ;
        RECT 15.330 20.465 15.500 20.635 ;
        RECT 15.330 20.105 15.500 20.275 ;
        RECT 15.330 19.745 15.500 19.915 ;
        RECT 15.330 19.385 15.500 19.555 ;
        RECT 15.330 19.025 15.500 19.195 ;
        RECT 15.330 18.665 15.500 18.835 ;
        RECT 15.330 18.305 15.500 18.475 ;
        RECT 15.330 17.945 15.500 18.115 ;
        RECT 15.330 17.585 15.500 17.755 ;
        RECT 15.330 17.225 15.500 17.395 ;
        RECT 15.330 16.865 15.500 17.035 ;
        RECT 15.330 16.505 15.500 16.675 ;
        RECT 15.330 16.145 15.500 16.315 ;
        RECT 15.330 15.785 15.500 15.955 ;
        RECT 16.910 21.185 17.080 21.355 ;
        RECT 16.910 20.825 17.080 20.995 ;
        RECT 16.910 20.465 17.080 20.635 ;
        RECT 16.910 20.105 17.080 20.275 ;
        RECT 16.910 19.745 17.080 19.915 ;
        RECT 16.910 19.385 17.080 19.555 ;
        RECT 16.910 19.025 17.080 19.195 ;
        RECT 16.910 18.665 17.080 18.835 ;
        RECT 16.910 18.305 17.080 18.475 ;
        RECT 16.910 17.945 17.080 18.115 ;
        RECT 16.910 17.585 17.080 17.755 ;
        RECT 16.910 17.225 17.080 17.395 ;
        RECT 16.910 16.865 17.080 17.035 ;
        RECT 16.910 16.505 17.080 16.675 ;
        RECT 16.910 16.145 17.080 16.315 ;
        RECT 16.910 15.785 17.080 15.955 ;
        RECT 18.490 21.185 18.660 21.355 ;
        RECT 18.490 20.825 18.660 20.995 ;
        RECT 18.490 20.465 18.660 20.635 ;
        RECT 28.740 20.365 28.910 20.535 ;
        RECT 29.100 20.365 29.270 20.535 ;
        RECT 29.460 20.365 29.630 20.535 ;
        RECT 29.820 20.365 29.990 20.535 ;
        RECT 30.180 20.365 30.350 20.535 ;
        RECT 30.540 20.365 30.710 20.535 ;
        RECT 30.900 20.365 31.070 20.535 ;
        RECT 31.260 20.365 31.430 20.535 ;
        RECT 31.620 20.365 31.790 20.535 ;
        RECT 31.980 20.365 32.150 20.535 ;
        RECT 32.340 20.365 32.510 20.535 ;
        RECT 32.700 20.365 32.870 20.535 ;
        RECT 33.060 20.365 33.230 20.535 ;
        RECT 33.420 20.365 33.590 20.535 ;
        RECT 33.780 20.365 33.950 20.535 ;
        RECT 34.140 20.365 34.310 20.535 ;
        RECT 34.500 20.365 34.670 20.535 ;
        RECT 34.860 20.365 35.030 20.535 ;
        RECT 35.220 20.365 35.390 20.535 ;
        RECT 35.580 20.365 35.750 20.535 ;
        RECT 35.940 20.365 36.110 20.535 ;
        RECT 36.300 20.365 36.470 20.535 ;
        RECT 36.660 20.365 36.830 20.535 ;
        RECT 37.020 20.365 37.190 20.535 ;
        RECT 37.380 20.365 37.550 20.535 ;
        RECT 37.740 20.365 37.910 20.535 ;
        RECT 38.100 20.365 38.270 20.535 ;
        RECT 38.460 20.365 38.630 20.535 ;
        RECT 38.820 20.365 38.990 20.535 ;
        RECT 39.180 20.365 39.350 20.535 ;
        RECT 39.540 20.365 39.710 20.535 ;
        RECT 39.900 20.365 40.070 20.535 ;
        RECT 40.260 20.365 40.430 20.535 ;
        RECT 40.620 20.365 40.790 20.535 ;
        RECT 40.980 20.365 41.150 20.535 ;
        RECT 41.340 20.365 41.510 20.535 ;
        RECT 41.700 20.365 41.870 20.535 ;
        RECT 42.060 20.365 42.230 20.535 ;
        RECT 42.420 20.365 42.590 20.535 ;
        RECT 42.780 20.365 42.950 20.535 ;
        RECT 43.140 20.365 43.310 20.535 ;
        RECT 43.500 20.365 43.670 20.535 ;
        RECT 43.860 20.365 44.030 20.535 ;
        RECT 44.220 20.365 44.390 20.535 ;
        RECT 44.580 20.365 44.750 20.535 ;
        RECT 44.940 20.365 45.110 20.535 ;
        RECT 45.300 20.365 45.470 20.535 ;
        RECT 45.660 20.365 45.830 20.535 ;
        RECT 46.020 20.365 46.190 20.535 ;
        RECT 46.380 20.365 46.550 20.535 ;
        RECT 46.740 20.365 46.910 20.535 ;
        RECT 47.100 20.365 47.270 20.535 ;
        RECT 47.460 20.365 47.630 20.535 ;
        RECT 18.490 20.105 18.660 20.275 ;
        RECT 18.490 19.745 18.660 19.915 ;
        RECT 18.490 19.385 18.660 19.555 ;
        RECT 18.490 19.025 18.660 19.195 ;
        RECT 18.490 18.665 18.660 18.835 ;
        RECT 18.490 18.305 18.660 18.475 ;
        RECT 18.490 17.945 18.660 18.115 ;
        RECT 18.490 17.585 18.660 17.755 ;
        RECT 18.490 17.225 18.660 17.395 ;
        RECT 18.490 16.865 18.660 17.035 ;
        RECT 18.490 16.505 18.660 16.675 ;
        RECT 18.490 16.145 18.660 16.315 ;
        RECT 18.490 15.785 18.660 15.955 ;
        RECT 3.165 14.990 3.335 15.160 ;
        RECT 3.525 14.990 3.695 15.160 ;
        RECT 3.885 14.990 4.055 15.160 ;
        RECT 4.245 14.990 4.415 15.160 ;
        RECT 4.605 14.990 4.775 15.160 ;
        RECT 4.965 14.990 5.135 15.160 ;
        RECT 5.325 14.990 5.495 15.160 ;
        RECT 5.685 14.990 5.855 15.160 ;
        RECT 6.045 14.990 6.215 15.160 ;
        RECT 6.405 14.990 6.575 15.160 ;
        RECT 6.765 14.990 6.935 15.160 ;
        RECT 7.125 14.990 7.295 15.160 ;
        RECT 7.485 14.990 7.655 15.160 ;
        RECT 7.845 14.990 8.015 15.160 ;
        RECT 8.205 14.990 8.375 15.160 ;
        RECT 8.565 14.990 8.735 15.160 ;
        RECT 8.925 14.990 9.095 15.160 ;
        RECT 9.285 14.990 9.455 15.160 ;
        RECT 9.645 14.990 9.815 15.160 ;
        RECT 10.005 14.990 10.175 15.160 ;
        RECT 10.365 14.990 10.535 15.160 ;
        RECT 10.725 14.990 10.895 15.160 ;
        RECT 11.085 14.990 11.255 15.160 ;
        RECT 11.445 14.990 11.615 15.160 ;
        RECT 11.805 14.990 11.975 15.160 ;
        RECT 12.165 14.990 12.335 15.160 ;
        RECT 12.525 14.990 12.695 15.160 ;
        RECT 12.885 14.990 13.055 15.160 ;
        RECT 13.245 14.990 13.415 15.160 ;
        RECT 13.605 14.990 13.775 15.160 ;
        RECT 13.965 14.990 14.135 15.160 ;
        RECT 14.325 14.990 14.495 15.160 ;
        RECT 14.685 14.990 14.855 15.160 ;
        RECT 15.045 14.990 15.215 15.160 ;
        RECT 15.405 14.990 15.575 15.160 ;
        RECT 15.765 14.990 15.935 15.160 ;
        RECT 16.125 14.990 16.295 15.160 ;
        RECT 16.485 14.990 16.655 15.160 ;
        RECT 16.845 14.990 17.015 15.160 ;
        RECT 17.205 14.990 17.375 15.160 ;
        RECT 17.565 14.990 17.735 15.160 ;
        RECT 17.925 14.990 18.095 15.160 ;
        RECT 2.370 8.390 2.540 8.560 ;
        RECT 2.370 8.030 2.540 8.200 ;
        RECT 2.370 7.670 2.540 7.840 ;
        RECT 2.370 7.310 2.540 7.480 ;
        RECT 2.370 6.950 2.540 7.120 ;
        RECT 2.370 6.590 2.540 6.760 ;
        RECT 2.370 6.230 2.540 6.400 ;
        RECT 2.370 5.870 2.540 6.040 ;
        RECT 2.370 5.510 2.540 5.680 ;
        RECT 2.370 5.150 2.540 5.320 ;
        RECT 2.370 4.790 2.540 4.960 ;
        RECT 2.370 4.430 2.540 4.600 ;
        RECT 2.370 4.070 2.540 4.240 ;
        RECT 2.370 3.710 2.540 3.880 ;
        RECT 3.160 8.390 3.330 8.560 ;
        RECT 3.160 8.030 3.330 8.200 ;
        RECT 3.160 7.670 3.330 7.840 ;
        RECT 3.160 7.310 3.330 7.480 ;
        RECT 3.160 6.950 3.330 7.120 ;
        RECT 3.160 6.590 3.330 6.760 ;
        RECT 3.160 6.230 3.330 6.400 ;
        RECT 3.160 5.870 3.330 6.040 ;
        RECT 3.160 5.510 3.330 5.680 ;
        RECT 3.160 5.150 3.330 5.320 ;
        RECT 3.160 4.790 3.330 4.960 ;
        RECT 3.160 4.430 3.330 4.600 ;
        RECT 3.160 4.070 3.330 4.240 ;
        RECT 3.160 3.710 3.330 3.880 ;
        RECT 3.950 8.390 4.120 8.560 ;
        RECT 3.950 8.030 4.120 8.200 ;
        RECT 3.950 7.670 4.120 7.840 ;
        RECT 3.950 7.310 4.120 7.480 ;
        RECT 3.950 6.950 4.120 7.120 ;
        RECT 3.950 6.590 4.120 6.760 ;
        RECT 3.950 6.230 4.120 6.400 ;
        RECT 3.950 5.870 4.120 6.040 ;
        RECT 3.950 5.510 4.120 5.680 ;
        RECT 3.950 5.150 4.120 5.320 ;
        RECT 3.950 4.790 4.120 4.960 ;
        RECT 3.950 4.430 4.120 4.600 ;
        RECT 3.950 4.070 4.120 4.240 ;
        RECT 3.950 3.710 4.120 3.880 ;
        RECT 4.740 8.390 4.910 8.560 ;
        RECT 4.740 8.030 4.910 8.200 ;
        RECT 4.740 7.670 4.910 7.840 ;
        RECT 4.740 7.310 4.910 7.480 ;
        RECT 4.740 6.950 4.910 7.120 ;
        RECT 4.740 6.590 4.910 6.760 ;
        RECT 4.740 6.230 4.910 6.400 ;
        RECT 4.740 5.870 4.910 6.040 ;
        RECT 4.740 5.510 4.910 5.680 ;
        RECT 4.740 5.150 4.910 5.320 ;
        RECT 4.740 4.790 4.910 4.960 ;
        RECT 4.740 4.430 4.910 4.600 ;
        RECT 4.740 4.070 4.910 4.240 ;
        RECT 4.740 3.710 4.910 3.880 ;
        RECT 5.530 8.390 5.700 8.560 ;
        RECT 5.530 8.030 5.700 8.200 ;
        RECT 5.530 7.670 5.700 7.840 ;
        RECT 5.530 7.310 5.700 7.480 ;
        RECT 5.530 6.950 5.700 7.120 ;
        RECT 5.530 6.590 5.700 6.760 ;
        RECT 5.530 6.230 5.700 6.400 ;
        RECT 5.530 5.870 5.700 6.040 ;
        RECT 5.530 5.510 5.700 5.680 ;
        RECT 5.530 5.150 5.700 5.320 ;
        RECT 5.530 4.790 5.700 4.960 ;
        RECT 5.530 4.430 5.700 4.600 ;
        RECT 5.530 4.070 5.700 4.240 ;
        RECT 5.530 3.710 5.700 3.880 ;
        RECT 6.320 8.390 6.490 8.560 ;
        RECT 6.320 8.030 6.490 8.200 ;
        RECT 6.320 7.670 6.490 7.840 ;
        RECT 6.320 7.310 6.490 7.480 ;
        RECT 6.320 6.950 6.490 7.120 ;
        RECT 6.320 6.590 6.490 6.760 ;
        RECT 6.320 6.230 6.490 6.400 ;
        RECT 6.320 5.870 6.490 6.040 ;
        RECT 6.320 5.510 6.490 5.680 ;
        RECT 6.320 5.150 6.490 5.320 ;
        RECT 6.320 4.790 6.490 4.960 ;
        RECT 6.320 4.430 6.490 4.600 ;
        RECT 6.320 4.070 6.490 4.240 ;
        RECT 6.320 3.710 6.490 3.880 ;
        RECT 7.110 8.390 7.280 8.560 ;
        RECT 7.110 8.030 7.280 8.200 ;
        RECT 7.110 7.670 7.280 7.840 ;
        RECT 7.110 7.310 7.280 7.480 ;
        RECT 7.110 6.950 7.280 7.120 ;
        RECT 7.110 6.590 7.280 6.760 ;
        RECT 7.110 6.230 7.280 6.400 ;
        RECT 7.110 5.870 7.280 6.040 ;
        RECT 7.110 5.510 7.280 5.680 ;
        RECT 7.110 5.150 7.280 5.320 ;
        RECT 7.110 4.790 7.280 4.960 ;
        RECT 7.110 4.430 7.280 4.600 ;
        RECT 7.110 4.070 7.280 4.240 ;
        RECT 7.110 3.710 7.280 3.880 ;
        RECT 7.900 8.390 8.070 8.560 ;
        RECT 7.900 8.030 8.070 8.200 ;
        RECT 7.900 7.670 8.070 7.840 ;
        RECT 7.900 7.310 8.070 7.480 ;
        RECT 7.900 6.950 8.070 7.120 ;
        RECT 7.900 6.590 8.070 6.760 ;
        RECT 7.900 6.230 8.070 6.400 ;
        RECT 7.900 5.870 8.070 6.040 ;
        RECT 7.900 5.510 8.070 5.680 ;
        RECT 7.900 5.150 8.070 5.320 ;
        RECT 7.900 4.790 8.070 4.960 ;
        RECT 7.900 4.430 8.070 4.600 ;
        RECT 7.900 4.070 8.070 4.240 ;
        RECT 7.900 3.710 8.070 3.880 ;
        RECT 8.690 8.390 8.860 8.560 ;
        RECT 8.690 8.030 8.860 8.200 ;
        RECT 8.690 7.670 8.860 7.840 ;
        RECT 8.690 7.310 8.860 7.480 ;
        RECT 8.690 6.950 8.860 7.120 ;
        RECT 8.690 6.590 8.860 6.760 ;
        RECT 8.690 6.230 8.860 6.400 ;
        RECT 8.690 5.870 8.860 6.040 ;
        RECT 8.690 5.510 8.860 5.680 ;
        RECT 8.690 5.150 8.860 5.320 ;
        RECT 8.690 4.790 8.860 4.960 ;
        RECT 8.690 4.430 8.860 4.600 ;
        RECT 8.690 4.070 8.860 4.240 ;
        RECT 8.690 3.710 8.860 3.880 ;
        RECT 9.480 8.390 9.650 8.560 ;
        RECT 9.480 8.030 9.650 8.200 ;
        RECT 9.480 7.670 9.650 7.840 ;
        RECT 9.480 7.310 9.650 7.480 ;
        RECT 9.480 6.950 9.650 7.120 ;
        RECT 9.480 6.590 9.650 6.760 ;
        RECT 9.480 6.230 9.650 6.400 ;
        RECT 9.480 5.870 9.650 6.040 ;
        RECT 9.480 5.510 9.650 5.680 ;
        RECT 9.480 5.150 9.650 5.320 ;
        RECT 9.480 4.790 9.650 4.960 ;
        RECT 9.480 4.430 9.650 4.600 ;
        RECT 9.480 4.070 9.650 4.240 ;
        RECT 9.480 3.710 9.650 3.880 ;
        RECT 10.270 8.390 10.440 8.560 ;
        RECT 10.270 8.030 10.440 8.200 ;
        RECT 10.270 7.670 10.440 7.840 ;
        RECT 10.270 7.310 10.440 7.480 ;
        RECT 10.270 6.950 10.440 7.120 ;
        RECT 10.270 6.590 10.440 6.760 ;
        RECT 10.270 6.230 10.440 6.400 ;
        RECT 10.270 5.870 10.440 6.040 ;
        RECT 10.270 5.510 10.440 5.680 ;
        RECT 10.270 5.150 10.440 5.320 ;
        RECT 10.270 4.790 10.440 4.960 ;
        RECT 10.270 4.430 10.440 4.600 ;
        RECT 10.270 4.070 10.440 4.240 ;
        RECT 10.270 3.710 10.440 3.880 ;
        RECT 11.060 8.390 11.230 8.560 ;
        RECT 11.060 8.030 11.230 8.200 ;
        RECT 11.060 7.670 11.230 7.840 ;
        RECT 11.060 7.310 11.230 7.480 ;
        RECT 11.060 6.950 11.230 7.120 ;
        RECT 11.060 6.590 11.230 6.760 ;
        RECT 11.060 6.230 11.230 6.400 ;
        RECT 11.060 5.870 11.230 6.040 ;
        RECT 11.060 5.510 11.230 5.680 ;
        RECT 11.060 5.150 11.230 5.320 ;
        RECT 11.060 4.790 11.230 4.960 ;
        RECT 11.060 4.430 11.230 4.600 ;
        RECT 11.060 4.070 11.230 4.240 ;
        RECT 11.060 3.710 11.230 3.880 ;
        RECT 11.850 8.390 12.020 8.560 ;
        RECT 11.850 8.030 12.020 8.200 ;
        RECT 11.850 7.670 12.020 7.840 ;
        RECT 11.850 7.310 12.020 7.480 ;
        RECT 11.850 6.950 12.020 7.120 ;
        RECT 11.850 6.590 12.020 6.760 ;
        RECT 11.850 6.230 12.020 6.400 ;
        RECT 11.850 5.870 12.020 6.040 ;
        RECT 11.850 5.510 12.020 5.680 ;
        RECT 11.850 5.150 12.020 5.320 ;
        RECT 11.850 4.790 12.020 4.960 ;
        RECT 11.850 4.430 12.020 4.600 ;
        RECT 11.850 4.070 12.020 4.240 ;
        RECT 11.850 3.710 12.020 3.880 ;
        RECT 12.640 8.390 12.810 8.560 ;
        RECT 12.640 8.030 12.810 8.200 ;
        RECT 12.640 7.670 12.810 7.840 ;
        RECT 12.640 7.310 12.810 7.480 ;
        RECT 12.640 6.950 12.810 7.120 ;
        RECT 12.640 6.590 12.810 6.760 ;
        RECT 12.640 6.230 12.810 6.400 ;
        RECT 12.640 5.870 12.810 6.040 ;
        RECT 12.640 5.510 12.810 5.680 ;
        RECT 12.640 5.150 12.810 5.320 ;
        RECT 12.640 4.790 12.810 4.960 ;
        RECT 12.640 4.430 12.810 4.600 ;
        RECT 12.640 4.070 12.810 4.240 ;
        RECT 12.640 3.710 12.810 3.880 ;
        RECT 13.430 8.390 13.600 8.560 ;
        RECT 13.430 8.030 13.600 8.200 ;
        RECT 13.430 7.670 13.600 7.840 ;
        RECT 13.430 7.310 13.600 7.480 ;
        RECT 13.430 6.950 13.600 7.120 ;
        RECT 13.430 6.590 13.600 6.760 ;
        RECT 13.430 6.230 13.600 6.400 ;
        RECT 13.430 5.870 13.600 6.040 ;
        RECT 13.430 5.510 13.600 5.680 ;
        RECT 13.430 5.150 13.600 5.320 ;
        RECT 13.430 4.790 13.600 4.960 ;
        RECT 13.430 4.430 13.600 4.600 ;
        RECT 13.430 4.070 13.600 4.240 ;
        RECT 13.430 3.710 13.600 3.880 ;
        RECT 14.220 8.390 14.390 8.560 ;
        RECT 14.220 8.030 14.390 8.200 ;
        RECT 14.220 7.670 14.390 7.840 ;
        RECT 14.220 7.310 14.390 7.480 ;
        RECT 14.220 6.950 14.390 7.120 ;
        RECT 14.220 6.590 14.390 6.760 ;
        RECT 14.220 6.230 14.390 6.400 ;
        RECT 14.220 5.870 14.390 6.040 ;
        RECT 14.220 5.510 14.390 5.680 ;
        RECT 14.220 5.150 14.390 5.320 ;
        RECT 14.220 4.790 14.390 4.960 ;
        RECT 14.220 4.430 14.390 4.600 ;
        RECT 14.220 4.070 14.390 4.240 ;
        RECT 14.220 3.710 14.390 3.880 ;
        RECT 15.010 8.390 15.180 8.560 ;
        RECT 15.010 8.030 15.180 8.200 ;
        RECT 15.010 7.670 15.180 7.840 ;
        RECT 15.010 7.310 15.180 7.480 ;
        RECT 15.010 6.950 15.180 7.120 ;
        RECT 15.010 6.590 15.180 6.760 ;
        RECT 15.010 6.230 15.180 6.400 ;
        RECT 15.010 5.870 15.180 6.040 ;
        RECT 15.010 5.510 15.180 5.680 ;
        RECT 15.010 5.150 15.180 5.320 ;
        RECT 15.010 4.790 15.180 4.960 ;
        RECT 15.010 4.430 15.180 4.600 ;
        RECT 15.010 4.070 15.180 4.240 ;
        RECT 15.010 3.710 15.180 3.880 ;
        RECT 15.800 8.390 15.970 8.560 ;
        RECT 15.800 8.030 15.970 8.200 ;
        RECT 15.800 7.670 15.970 7.840 ;
        RECT 15.800 7.310 15.970 7.480 ;
        RECT 15.800 6.950 15.970 7.120 ;
        RECT 15.800 6.590 15.970 6.760 ;
        RECT 15.800 6.230 15.970 6.400 ;
        RECT 15.800 5.870 15.970 6.040 ;
        RECT 15.800 5.510 15.970 5.680 ;
        RECT 15.800 5.150 15.970 5.320 ;
        RECT 15.800 4.790 15.970 4.960 ;
        RECT 15.800 4.430 15.970 4.600 ;
        RECT 15.800 4.070 15.970 4.240 ;
        RECT 15.800 3.710 15.970 3.880 ;
        RECT 16.590 8.390 16.760 8.560 ;
        RECT 16.590 8.030 16.760 8.200 ;
        RECT 16.590 7.670 16.760 7.840 ;
        RECT 16.590 7.310 16.760 7.480 ;
        RECT 16.590 6.950 16.760 7.120 ;
        RECT 16.590 6.590 16.760 6.760 ;
        RECT 16.590 6.230 16.760 6.400 ;
        RECT 16.590 5.870 16.760 6.040 ;
        RECT 16.590 5.510 16.760 5.680 ;
        RECT 16.590 5.150 16.760 5.320 ;
        RECT 16.590 4.790 16.760 4.960 ;
        RECT 16.590 4.430 16.760 4.600 ;
        RECT 16.590 4.070 16.760 4.240 ;
        RECT 16.590 3.710 16.760 3.880 ;
        RECT 17.380 8.390 17.550 8.560 ;
        RECT 17.380 8.030 17.550 8.200 ;
        RECT 17.380 7.670 17.550 7.840 ;
        RECT 17.380 7.310 17.550 7.480 ;
        RECT 17.380 6.950 17.550 7.120 ;
        RECT 17.380 6.590 17.550 6.760 ;
        RECT 17.380 6.230 17.550 6.400 ;
        RECT 17.380 5.870 17.550 6.040 ;
        RECT 17.380 5.510 17.550 5.680 ;
        RECT 17.380 5.150 17.550 5.320 ;
        RECT 17.380 4.790 17.550 4.960 ;
        RECT 17.380 4.430 17.550 4.600 ;
        RECT 17.380 4.070 17.550 4.240 ;
        RECT 17.380 3.710 17.550 3.880 ;
        RECT 18.170 8.390 18.340 8.560 ;
        RECT 18.170 8.030 18.340 8.200 ;
        RECT 18.170 7.670 18.340 7.840 ;
        RECT 18.170 7.310 18.340 7.480 ;
        RECT 18.170 6.950 18.340 7.120 ;
        RECT 18.170 6.590 18.340 6.760 ;
        RECT 18.170 6.230 18.340 6.400 ;
        RECT 18.170 5.870 18.340 6.040 ;
        RECT 18.170 5.510 18.340 5.680 ;
        RECT 18.170 5.150 18.340 5.320 ;
        RECT 28.740 5.165 28.910 5.335 ;
        RECT 29.100 5.165 29.270 5.335 ;
        RECT 29.460 5.165 29.630 5.335 ;
        RECT 29.820 5.165 29.990 5.335 ;
        RECT 30.180 5.165 30.350 5.335 ;
        RECT 30.540 5.165 30.710 5.335 ;
        RECT 30.900 5.165 31.070 5.335 ;
        RECT 31.260 5.165 31.430 5.335 ;
        RECT 31.620 5.165 31.790 5.335 ;
        RECT 31.980 5.165 32.150 5.335 ;
        RECT 32.340 5.165 32.510 5.335 ;
        RECT 32.700 5.165 32.870 5.335 ;
        RECT 33.060 5.165 33.230 5.335 ;
        RECT 33.420 5.165 33.590 5.335 ;
        RECT 33.780 5.165 33.950 5.335 ;
        RECT 34.140 5.165 34.310 5.335 ;
        RECT 34.500 5.165 34.670 5.335 ;
        RECT 34.860 5.165 35.030 5.335 ;
        RECT 35.220 5.165 35.390 5.335 ;
        RECT 35.580 5.165 35.750 5.335 ;
        RECT 35.940 5.165 36.110 5.335 ;
        RECT 36.300 5.165 36.470 5.335 ;
        RECT 36.660 5.165 36.830 5.335 ;
        RECT 37.020 5.165 37.190 5.335 ;
        RECT 37.380 5.165 37.550 5.335 ;
        RECT 37.740 5.165 37.910 5.335 ;
        RECT 38.100 5.165 38.270 5.335 ;
        RECT 38.460 5.165 38.630 5.335 ;
        RECT 38.820 5.165 38.990 5.335 ;
        RECT 39.180 5.165 39.350 5.335 ;
        RECT 39.540 5.165 39.710 5.335 ;
        RECT 39.900 5.165 40.070 5.335 ;
        RECT 40.260 5.165 40.430 5.335 ;
        RECT 40.620 5.165 40.790 5.335 ;
        RECT 40.980 5.165 41.150 5.335 ;
        RECT 41.340 5.165 41.510 5.335 ;
        RECT 41.700 5.165 41.870 5.335 ;
        RECT 42.060 5.165 42.230 5.335 ;
        RECT 42.420 5.165 42.590 5.335 ;
        RECT 42.780 5.165 42.950 5.335 ;
        RECT 43.140 5.165 43.310 5.335 ;
        RECT 43.500 5.165 43.670 5.335 ;
        RECT 43.860 5.165 44.030 5.335 ;
        RECT 44.220 5.165 44.390 5.335 ;
        RECT 44.580 5.165 44.750 5.335 ;
        RECT 44.940 5.165 45.110 5.335 ;
        RECT 45.300 5.165 45.470 5.335 ;
        RECT 45.660 5.165 45.830 5.335 ;
        RECT 46.020 5.165 46.190 5.335 ;
        RECT 46.380 5.165 46.550 5.335 ;
        RECT 46.740 5.165 46.910 5.335 ;
        RECT 47.100 5.165 47.270 5.335 ;
        RECT 47.460 5.165 47.630 5.335 ;
        RECT 18.170 4.790 18.340 4.960 ;
        RECT 18.170 4.430 18.340 4.600 ;
        RECT 18.170 4.070 18.340 4.240 ;
        RECT 18.170 3.710 18.340 3.880 ;
        RECT 4.810 -2.190 4.980 -2.020 ;
        RECT 4.810 -2.550 4.980 -2.380 ;
        RECT 4.810 -2.910 4.980 -2.740 ;
        RECT 4.810 -3.270 4.980 -3.100 ;
        RECT 4.810 -3.630 4.980 -3.460 ;
        RECT 4.810 -3.990 4.980 -3.820 ;
        RECT 4.810 -4.350 4.980 -4.180 ;
        RECT 4.810 -4.710 4.980 -4.540 ;
        RECT 4.810 -5.070 4.980 -4.900 ;
        RECT 4.810 -5.430 4.980 -5.260 ;
        RECT 4.810 -5.790 4.980 -5.620 ;
        RECT 4.810 -6.150 4.980 -5.980 ;
        RECT 4.810 -6.510 4.980 -6.340 ;
        RECT 4.810 -6.870 4.980 -6.700 ;
        RECT 4.810 -7.230 4.980 -7.060 ;
        RECT 4.810 -7.590 4.980 -7.420 ;
        RECT 4.810 -7.950 4.980 -7.780 ;
        RECT 4.810 -8.310 4.980 -8.140 ;
        RECT 4.810 -8.670 4.980 -8.500 ;
        RECT 4.810 -9.030 4.980 -8.860 ;
        RECT 4.810 -9.390 4.980 -9.220 ;
        RECT 4.810 -9.750 4.980 -9.580 ;
        RECT 4.810 -10.110 4.980 -9.940 ;
        RECT 4.810 -10.470 4.980 -10.300 ;
        RECT 4.810 -10.830 4.980 -10.660 ;
        RECT 4.810 -11.190 4.980 -11.020 ;
        RECT 4.810 -11.550 4.980 -11.380 ;
        RECT 4.810 -11.910 4.980 -11.740 ;
        RECT 4.810 -12.270 4.980 -12.100 ;
      LAYER met1 ;
        RECT 2.065 21.910 19.365 22.230 ;
        RECT 2.065 16.300 2.440 21.910 ;
        RECT 2.660 16.300 2.890 21.570 ;
        RECT 4.240 21.355 4.470 21.570 ;
        RECT 4.195 20.775 4.515 21.355 ;
        RECT 2.065 15.720 2.935 16.300 ;
        RECT 2.065 15.230 2.440 15.720 ;
        RECT 2.660 15.570 2.890 15.720 ;
        RECT 4.240 15.570 4.470 20.775 ;
        RECT 5.820 16.300 6.050 21.570 ;
        RECT 7.400 21.355 7.630 21.570 ;
        RECT 7.355 20.775 7.675 21.355 ;
        RECT 5.775 15.720 6.095 16.300 ;
        RECT 5.820 15.570 6.050 15.720 ;
        RECT 7.400 15.570 7.630 20.775 ;
        RECT 8.980 16.300 9.210 21.570 ;
        RECT 10.560 21.355 10.790 21.570 ;
        RECT 10.515 20.775 10.835 21.355 ;
        RECT 8.935 15.720 9.255 16.300 ;
        RECT 8.980 15.570 9.210 15.720 ;
        RECT 10.560 15.570 10.790 20.775 ;
        RECT 12.140 16.300 12.370 21.570 ;
        RECT 13.720 21.355 13.950 21.570 ;
        RECT 13.675 20.775 13.995 21.355 ;
        RECT 12.095 15.720 12.415 16.300 ;
        RECT 12.140 15.570 12.370 15.720 ;
        RECT 13.720 15.570 13.950 20.775 ;
        RECT 15.300 16.300 15.530 21.570 ;
        RECT 16.880 21.355 17.110 21.570 ;
        RECT 16.835 20.775 17.155 21.355 ;
        RECT 15.255 15.720 15.575 16.300 ;
        RECT 15.300 15.570 15.530 15.720 ;
        RECT 16.880 15.570 17.110 20.775 ;
        RECT 18.460 16.300 18.690 21.570 ;
        RECT 18.990 16.300 19.365 21.910 ;
        RECT 18.415 15.720 19.365 16.300 ;
        RECT 18.460 15.570 18.690 15.720 ;
        RECT 18.990 15.230 19.365 15.720 ;
        RECT 2.065 14.910 19.365 15.230 ;
        RECT 27.020 20.605 27.870 21.355 ;
        RECT 27.020 20.285 49.350 20.605 ;
        RECT 2.340 4.445 2.570 8.635 ;
        RECT 3.130 6.600 3.360 8.635 ;
        RECT 3.920 8.300 4.150 8.635 ;
        RECT 3.875 7.735 4.195 8.300 ;
        RECT 3.100 6.020 3.390 6.600 ;
        RECT 2.295 3.875 2.615 4.445 ;
        RECT 2.340 3.635 2.570 3.875 ;
        RECT 3.130 3.635 3.360 6.020 ;
        RECT 3.920 3.635 4.150 7.735 ;
        RECT 4.710 6.600 4.940 8.635 ;
        RECT 4.680 6.020 4.970 6.600 ;
        RECT 4.710 3.635 4.940 6.020 ;
        RECT 5.500 4.445 5.730 8.635 ;
        RECT 6.290 6.600 6.520 8.635 ;
        RECT 7.080 8.300 7.310 8.635 ;
        RECT 7.035 7.735 7.355 8.300 ;
        RECT 6.260 6.020 6.550 6.600 ;
        RECT 5.455 3.875 5.775 4.445 ;
        RECT 5.500 3.635 5.730 3.875 ;
        RECT 6.290 3.635 6.520 6.020 ;
        RECT 7.080 3.635 7.310 7.735 ;
        RECT 7.870 6.600 8.100 8.635 ;
        RECT 7.840 6.020 8.130 6.600 ;
        RECT 7.870 3.635 8.100 6.020 ;
        RECT 8.660 4.445 8.890 8.635 ;
        RECT 9.450 6.600 9.680 8.635 ;
        RECT 10.240 8.300 10.470 8.635 ;
        RECT 10.195 7.735 10.515 8.300 ;
        RECT 9.420 6.020 9.710 6.600 ;
        RECT 8.615 3.875 8.935 4.445 ;
        RECT 8.660 3.635 8.890 3.875 ;
        RECT 9.450 3.635 9.680 6.020 ;
        RECT 10.240 3.635 10.470 7.735 ;
        RECT 11.030 6.600 11.260 8.635 ;
        RECT 11.000 6.020 11.290 6.600 ;
        RECT 11.030 3.635 11.260 6.020 ;
        RECT 11.820 4.445 12.050 8.635 ;
        RECT 12.610 6.600 12.840 8.635 ;
        RECT 13.400 8.300 13.630 8.635 ;
        RECT 13.355 7.735 13.675 8.300 ;
        RECT 12.580 6.020 12.870 6.600 ;
        RECT 11.775 3.875 12.095 4.445 ;
        RECT 11.820 3.635 12.050 3.875 ;
        RECT 12.610 3.635 12.840 6.020 ;
        RECT 13.400 3.635 13.630 7.735 ;
        RECT 14.190 6.600 14.420 8.635 ;
        RECT 14.160 6.020 14.450 6.600 ;
        RECT 14.190 3.635 14.420 6.020 ;
        RECT 14.980 4.445 15.210 8.635 ;
        RECT 15.770 6.600 16.000 8.635 ;
        RECT 16.560 8.300 16.790 8.635 ;
        RECT 16.515 7.735 16.835 8.300 ;
        RECT 15.740 6.020 16.030 6.600 ;
        RECT 14.935 3.875 15.255 4.445 ;
        RECT 14.980 3.635 15.210 3.875 ;
        RECT 15.770 3.635 16.000 6.020 ;
        RECT 16.560 3.635 16.790 7.735 ;
        RECT 17.350 6.600 17.580 8.635 ;
        RECT 17.320 6.020 17.610 6.600 ;
        RECT 17.350 3.635 17.580 6.020 ;
        RECT 18.140 4.445 18.370 8.635 ;
        RECT 27.020 5.405 27.870 20.285 ;
        RECT 48.500 5.405 49.350 20.285 ;
        RECT 27.020 5.085 49.350 5.405 ;
        RECT 18.095 3.875 18.415 4.445 ;
        RECT 18.140 3.635 18.370 3.875 ;
        RECT 4.780 -3.675 5.010 -1.895 ;
        RECT 4.735 -4.725 5.055 -3.675 ;
        RECT 4.780 -12.395 5.010 -4.725 ;
      LAYER via ;
        RECT 4.225 20.935 4.485 21.195 ;
        RECT 2.645 15.880 2.905 16.140 ;
        RECT 7.385 20.935 7.645 21.195 ;
        RECT 5.805 15.880 6.065 16.140 ;
        RECT 10.545 20.935 10.805 21.195 ;
        RECT 8.965 15.880 9.225 16.140 ;
        RECT 13.705 20.935 13.965 21.195 ;
        RECT 12.125 15.880 12.385 16.140 ;
        RECT 16.865 20.935 17.125 21.195 ;
        RECT 15.285 15.880 15.545 16.140 ;
        RECT 18.445 15.880 18.705 16.140 ;
        RECT 27.155 20.555 27.735 21.135 ;
        RECT 3.905 7.885 4.165 8.145 ;
        RECT 3.115 6.170 3.375 6.430 ;
        RECT 2.325 4.025 2.585 4.285 ;
        RECT 4.695 6.170 4.955 6.430 ;
        RECT 7.065 7.885 7.325 8.145 ;
        RECT 6.275 6.170 6.535 6.430 ;
        RECT 5.485 4.025 5.745 4.285 ;
        RECT 7.855 6.170 8.115 6.430 ;
        RECT 10.225 7.885 10.485 8.145 ;
        RECT 9.435 6.170 9.695 6.430 ;
        RECT 8.645 4.025 8.905 4.285 ;
        RECT 11.015 6.170 11.275 6.430 ;
        RECT 13.385 7.885 13.645 8.145 ;
        RECT 12.595 6.170 12.855 6.430 ;
        RECT 11.805 4.025 12.065 4.285 ;
        RECT 14.175 6.170 14.435 6.430 ;
        RECT 16.545 7.885 16.805 8.145 ;
        RECT 15.755 6.170 16.015 6.430 ;
        RECT 14.965 4.025 15.225 4.285 ;
        RECT 17.335 6.170 17.595 6.430 ;
        RECT 18.125 4.025 18.385 4.285 ;
        RECT 4.765 -4.010 5.025 -3.750 ;
        RECT 4.765 -4.330 5.025 -4.070 ;
        RECT 4.765 -4.650 5.025 -4.390 ;
      LAYER met2 ;
        RECT -0.090 20.775 27.870 21.355 ;
        RECT 27.020 20.275 27.870 20.775 ;
        RECT 2.630 15.720 18.720 16.300 ;
        RECT 2.310 7.735 18.400 8.315 ;
        RECT 2.310 6.020 18.400 6.600 ;
        RECT 2.310 3.875 18.400 4.455 ;
        RECT 3.170 -4.745 11.360 -3.665 ;
      LAYER via2 ;
        RECT 5.125 20.915 5.405 21.195 ;
        RECT 13.025 20.930 13.305 21.210 ;
        RECT 20.735 20.910 21.015 21.190 ;
        RECT 21.135 20.910 21.415 21.190 ;
        RECT 21.535 20.910 21.815 21.190 ;
        RECT 21.935 20.910 22.215 21.190 ;
        RECT 22.335 20.910 22.615 21.190 ;
        RECT 22.735 20.910 23.015 21.190 ;
        RECT 23.135 20.910 23.415 21.190 ;
        RECT 23.535 20.910 23.815 21.190 ;
        RECT 3.025 15.845 3.305 16.125 ;
        RECT 18.015 15.865 18.295 16.145 ;
        RECT 5.095 7.885 5.375 8.165 ;
        RECT 12.990 7.880 13.270 8.160 ;
        RECT 4.505 6.165 4.785 6.445 ;
        RECT 4.905 6.165 5.185 6.445 ;
        RECT 7.665 6.170 7.945 6.450 ;
        RECT 8.065 6.170 8.345 6.450 ;
        RECT 2.710 4.040 2.990 4.320 ;
        RECT 17.715 4.040 17.995 4.320 ;
        RECT 4.500 -4.560 5.180 -3.880 ;
        RECT 7.680 -4.555 8.360 -3.875 ;
      LAYER met3 ;
        RECT 2.295 3.875 3.475 16.300 ;
        RECT 4.940 7.735 5.600 21.355 ;
        RECT 12.840 7.735 13.500 21.355 ;
        RECT 4.220 -4.745 5.470 6.600 ;
        RECT 7.380 -4.745 8.630 6.600 ;
        RECT 17.255 3.875 18.435 16.300 ;
        RECT 20.585 -15.085 23.985 21.355 ;
      LAYER via3 ;
        RECT 20.900 -14.725 23.620 -4.005 ;
      LAYER met4 ;
        RECT 28.320 -3.370 51.930 -0.330 ;
        RECT 20.585 -15.085 51.930 -3.370 ;
        RECT 28.320 -23.940 51.930 -15.085 ;
  END
END OpampM
END LIBRARY

