magic
tech sky130A
magscale 1 2
timestamp 1667243390
<< obsli1 >>
rect 1104 2159 248860 247537
<< obsm1 >>
rect 14 1776 248860 247568
<< metal2 >>
rect 662 249200 718 250000
rect 1950 249200 2006 250000
rect 3882 249200 3938 250000
rect 5170 249200 5226 250000
rect 7102 249200 7158 250000
rect 8390 249200 8446 250000
rect 10322 249200 10378 250000
rect 11610 249200 11666 250000
rect 13542 249200 13598 250000
rect 14830 249200 14886 250000
rect 16762 249200 16818 250000
rect 18050 249200 18106 250000
rect 19982 249200 20038 250000
rect 21270 249200 21326 250000
rect 23202 249200 23258 250000
rect 24490 249200 24546 250000
rect 26422 249200 26478 250000
rect 27710 249200 27766 250000
rect 29642 249200 29698 250000
rect 30930 249200 30986 250000
rect 32862 249200 32918 250000
rect 34150 249200 34206 250000
rect 36082 249200 36138 250000
rect 37370 249200 37426 250000
rect 39302 249200 39358 250000
rect 40590 249200 40646 250000
rect 41878 249200 41934 250000
rect 43810 249200 43866 250000
rect 45098 249200 45154 250000
rect 47030 249200 47086 250000
rect 48318 249200 48374 250000
rect 50250 249200 50306 250000
rect 51538 249200 51594 250000
rect 53470 249200 53526 250000
rect 54758 249200 54814 250000
rect 56690 249200 56746 250000
rect 57978 249200 58034 250000
rect 59910 249200 59966 250000
rect 61198 249200 61254 250000
rect 63130 249200 63186 250000
rect 64418 249200 64474 250000
rect 66350 249200 66406 250000
rect 67638 249200 67694 250000
rect 69570 249200 69626 250000
rect 70858 249200 70914 250000
rect 72790 249200 72846 250000
rect 74078 249200 74134 250000
rect 76010 249200 76066 250000
rect 77298 249200 77354 250000
rect 79230 249200 79286 250000
rect 80518 249200 80574 250000
rect 82450 249200 82506 250000
rect 83738 249200 83794 250000
rect 85670 249200 85726 250000
rect 86958 249200 87014 250000
rect 88890 249200 88946 250000
rect 90178 249200 90234 250000
rect 92110 249200 92166 250000
rect 93398 249200 93454 250000
rect 95330 249200 95386 250000
rect 96618 249200 96674 250000
rect 98550 249200 98606 250000
rect 99838 249200 99894 250000
rect 101770 249200 101826 250000
rect 103058 249200 103114 250000
rect 104990 249200 105046 250000
rect 106278 249200 106334 250000
rect 108210 249200 108266 250000
rect 109498 249200 109554 250000
rect 111430 249200 111486 250000
rect 112718 249200 112774 250000
rect 114650 249200 114706 250000
rect 115938 249200 115994 250000
rect 117870 249200 117926 250000
rect 119158 249200 119214 250000
rect 121090 249200 121146 250000
rect 122378 249200 122434 250000
rect 124310 249200 124366 250000
rect 125598 249200 125654 250000
rect 127530 249200 127586 250000
rect 128818 249200 128874 250000
rect 130750 249200 130806 250000
rect 132038 249200 132094 250000
rect 133970 249200 134026 250000
rect 135258 249200 135314 250000
rect 137190 249200 137246 250000
rect 138478 249200 138534 250000
rect 140410 249200 140466 250000
rect 141698 249200 141754 250000
rect 143630 249200 143686 250000
rect 144918 249200 144974 250000
rect 146850 249200 146906 250000
rect 148138 249200 148194 250000
rect 150070 249200 150126 250000
rect 151358 249200 151414 250000
rect 153290 249200 153346 250000
rect 154578 249200 154634 250000
rect 156510 249200 156566 250000
rect 157798 249200 157854 250000
rect 159730 249200 159786 250000
rect 161018 249200 161074 250000
rect 162950 249200 163006 250000
rect 164238 249200 164294 250000
rect 166170 249200 166226 250000
rect 167458 249200 167514 250000
rect 169390 249200 169446 250000
rect 170678 249200 170734 250000
rect 172610 249200 172666 250000
rect 173898 249200 173954 250000
rect 175830 249200 175886 250000
rect 177118 249200 177174 250000
rect 179050 249200 179106 250000
rect 180338 249200 180394 250000
rect 181626 249200 181682 250000
rect 183558 249200 183614 250000
rect 184846 249200 184902 250000
rect 186778 249200 186834 250000
rect 188066 249200 188122 250000
rect 189998 249200 190054 250000
rect 191286 249200 191342 250000
rect 193218 249200 193274 250000
rect 194506 249200 194562 250000
rect 196438 249200 196494 250000
rect 197726 249200 197782 250000
rect 199658 249200 199714 250000
rect 200946 249200 201002 250000
rect 202878 249200 202934 250000
rect 204166 249200 204222 250000
rect 206098 249200 206154 250000
rect 207386 249200 207442 250000
rect 209318 249200 209374 250000
rect 210606 249200 210662 250000
rect 212538 249200 212594 250000
rect 213826 249200 213882 250000
rect 215758 249200 215814 250000
rect 217046 249200 217102 250000
rect 218978 249200 219034 250000
rect 220266 249200 220322 250000
rect 222198 249200 222254 250000
rect 223486 249200 223542 250000
rect 225418 249200 225474 250000
rect 226706 249200 226762 250000
rect 228638 249200 228694 250000
rect 229926 249200 229982 250000
rect 231858 249200 231914 250000
rect 233146 249200 233202 250000
rect 235078 249200 235134 250000
rect 236366 249200 236422 250000
rect 238298 249200 238354 250000
rect 239586 249200 239642 250000
rect 241518 249200 241574 250000
rect 242806 249200 242862 250000
rect 244738 249200 244794 250000
rect 246026 249200 246082 250000
rect 247958 249200 248014 250000
rect 249246 249200 249302 250000
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36726 0 36782 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 43166 0 43222 800
rect 44454 0 44510 800
rect 46386 0 46442 800
rect 47674 0 47730 800
rect 49606 0 49662 800
rect 50894 0 50950 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 59266 0 59322 800
rect 60554 0 60610 800
rect 62486 0 62542 800
rect 63774 0 63830 800
rect 65706 0 65762 800
rect 66994 0 67050 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 72146 0 72202 800
rect 73434 0 73490 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 78586 0 78642 800
rect 79874 0 79930 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 85026 0 85082 800
rect 86314 0 86370 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 91466 0 91522 800
rect 92754 0 92810 800
rect 94686 0 94742 800
rect 95974 0 96030 800
rect 97906 0 97962 800
rect 99194 0 99250 800
rect 101126 0 101182 800
rect 102414 0 102470 800
rect 104346 0 104402 800
rect 105634 0 105690 800
rect 107566 0 107622 800
rect 108854 0 108910 800
rect 110786 0 110842 800
rect 112074 0 112130 800
rect 114006 0 114062 800
rect 115294 0 115350 800
rect 117226 0 117282 800
rect 118514 0 118570 800
rect 120446 0 120502 800
rect 121734 0 121790 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 126886 0 126942 800
rect 128174 0 128230 800
rect 130106 0 130162 800
rect 131394 0 131450 800
rect 133326 0 133382 800
rect 134614 0 134670 800
rect 136546 0 136602 800
rect 137834 0 137890 800
rect 139122 0 139178 800
rect 141054 0 141110 800
rect 142342 0 142398 800
rect 144274 0 144330 800
rect 145562 0 145618 800
rect 147494 0 147550 800
rect 148782 0 148838 800
rect 150714 0 150770 800
rect 152002 0 152058 800
rect 153934 0 153990 800
rect 155222 0 155278 800
rect 157154 0 157210 800
rect 158442 0 158498 800
rect 160374 0 160430 800
rect 161662 0 161718 800
rect 163594 0 163650 800
rect 164882 0 164938 800
rect 166814 0 166870 800
rect 168102 0 168158 800
rect 170034 0 170090 800
rect 171322 0 171378 800
rect 173254 0 173310 800
rect 174542 0 174598 800
rect 176474 0 176530 800
rect 177762 0 177818 800
rect 179694 0 179750 800
rect 180982 0 181038 800
rect 182914 0 182970 800
rect 184202 0 184258 800
rect 186134 0 186190 800
rect 187422 0 187478 800
rect 189354 0 189410 800
rect 190642 0 190698 800
rect 192574 0 192630 800
rect 193862 0 193918 800
rect 195794 0 195850 800
rect 197082 0 197138 800
rect 199014 0 199070 800
rect 200302 0 200358 800
rect 202234 0 202290 800
rect 203522 0 203578 800
rect 205454 0 205510 800
rect 206742 0 206798 800
rect 208674 0 208730 800
rect 209962 0 210018 800
rect 211894 0 211950 800
rect 213182 0 213238 800
rect 215114 0 215170 800
rect 216402 0 216458 800
rect 218334 0 218390 800
rect 219622 0 219678 800
rect 221554 0 221610 800
rect 222842 0 222898 800
rect 224774 0 224830 800
rect 226062 0 226118 800
rect 227994 0 228050 800
rect 229282 0 229338 800
rect 231214 0 231270 800
rect 232502 0 232558 800
rect 234434 0 234490 800
rect 235722 0 235778 800
rect 237654 0 237710 800
rect 238942 0 238998 800
rect 240874 0 240930 800
rect 242162 0 242218 800
rect 244094 0 244150 800
rect 245382 0 245438 800
rect 247314 0 247370 800
rect 248602 0 248658 800
<< obsm2 >>
rect 20 249144 606 249234
rect 774 249144 1894 249234
rect 2062 249144 3826 249234
rect 3994 249144 5114 249234
rect 5282 249144 7046 249234
rect 7214 249144 8334 249234
rect 8502 249144 10266 249234
rect 10434 249144 11554 249234
rect 11722 249144 13486 249234
rect 13654 249144 14774 249234
rect 14942 249144 16706 249234
rect 16874 249144 17994 249234
rect 18162 249144 19926 249234
rect 20094 249144 21214 249234
rect 21382 249144 23146 249234
rect 23314 249144 24434 249234
rect 24602 249144 26366 249234
rect 26534 249144 27654 249234
rect 27822 249144 29586 249234
rect 29754 249144 30874 249234
rect 31042 249144 32806 249234
rect 32974 249144 34094 249234
rect 34262 249144 36026 249234
rect 36194 249144 37314 249234
rect 37482 249144 39246 249234
rect 39414 249144 40534 249234
rect 40702 249144 41822 249234
rect 41990 249144 43754 249234
rect 43922 249144 45042 249234
rect 45210 249144 46974 249234
rect 47142 249144 48262 249234
rect 48430 249144 50194 249234
rect 50362 249144 51482 249234
rect 51650 249144 53414 249234
rect 53582 249144 54702 249234
rect 54870 249144 56634 249234
rect 56802 249144 57922 249234
rect 58090 249144 59854 249234
rect 60022 249144 61142 249234
rect 61310 249144 63074 249234
rect 63242 249144 64362 249234
rect 64530 249144 66294 249234
rect 66462 249144 67582 249234
rect 67750 249144 69514 249234
rect 69682 249144 70802 249234
rect 70970 249144 72734 249234
rect 72902 249144 74022 249234
rect 74190 249144 75954 249234
rect 76122 249144 77242 249234
rect 77410 249144 79174 249234
rect 79342 249144 80462 249234
rect 80630 249144 82394 249234
rect 82562 249144 83682 249234
rect 83850 249144 85614 249234
rect 85782 249144 86902 249234
rect 87070 249144 88834 249234
rect 89002 249144 90122 249234
rect 90290 249144 92054 249234
rect 92222 249144 93342 249234
rect 93510 249144 95274 249234
rect 95442 249144 96562 249234
rect 96730 249144 98494 249234
rect 98662 249144 99782 249234
rect 99950 249144 101714 249234
rect 101882 249144 103002 249234
rect 103170 249144 104934 249234
rect 105102 249144 106222 249234
rect 106390 249144 108154 249234
rect 108322 249144 109442 249234
rect 109610 249144 111374 249234
rect 111542 249144 112662 249234
rect 112830 249144 114594 249234
rect 114762 249144 115882 249234
rect 116050 249144 117814 249234
rect 117982 249144 119102 249234
rect 119270 249144 121034 249234
rect 121202 249144 122322 249234
rect 122490 249144 124254 249234
rect 124422 249144 125542 249234
rect 125710 249144 127474 249234
rect 127642 249144 128762 249234
rect 128930 249144 130694 249234
rect 130862 249144 131982 249234
rect 132150 249144 133914 249234
rect 134082 249144 135202 249234
rect 135370 249144 137134 249234
rect 137302 249144 138422 249234
rect 138590 249144 140354 249234
rect 140522 249144 141642 249234
rect 141810 249144 143574 249234
rect 143742 249144 144862 249234
rect 145030 249144 146794 249234
rect 146962 249144 148082 249234
rect 148250 249144 150014 249234
rect 150182 249144 151302 249234
rect 151470 249144 153234 249234
rect 153402 249144 154522 249234
rect 154690 249144 156454 249234
rect 156622 249144 157742 249234
rect 157910 249144 159674 249234
rect 159842 249144 160962 249234
rect 161130 249144 162894 249234
rect 163062 249144 164182 249234
rect 164350 249144 166114 249234
rect 166282 249144 167402 249234
rect 167570 249144 169334 249234
rect 169502 249144 170622 249234
rect 170790 249144 172554 249234
rect 172722 249144 173842 249234
rect 174010 249144 175774 249234
rect 175942 249144 177062 249234
rect 177230 249144 178994 249234
rect 179162 249144 180282 249234
rect 180450 249144 181570 249234
rect 181738 249144 183502 249234
rect 183670 249144 184790 249234
rect 184958 249144 186722 249234
rect 186890 249144 188010 249234
rect 188178 249144 189942 249234
rect 190110 249144 191230 249234
rect 191398 249144 193162 249234
rect 193330 249144 194450 249234
rect 194618 249144 196382 249234
rect 196550 249144 197670 249234
rect 197838 249144 199602 249234
rect 199770 249144 200890 249234
rect 201058 249144 202822 249234
rect 202990 249144 204110 249234
rect 204278 249144 206042 249234
rect 206210 249144 207330 249234
rect 207498 249144 209262 249234
rect 209430 249144 210550 249234
rect 210718 249144 212482 249234
rect 212650 249144 213770 249234
rect 213938 249144 215702 249234
rect 215870 249144 216990 249234
rect 217158 249144 218922 249234
rect 219090 249144 220210 249234
rect 220378 249144 222142 249234
rect 222310 249144 223430 249234
rect 223598 249144 225362 249234
rect 225530 249144 226650 249234
rect 226818 249144 228582 249234
rect 228750 249144 229870 249234
rect 230038 249144 231802 249234
rect 231970 249144 233090 249234
rect 233258 249144 235022 249234
rect 235190 249144 236310 249234
rect 236478 249144 238242 249234
rect 238410 249144 239530 249234
rect 239698 249144 241462 249234
rect 241630 249144 242750 249234
rect 242918 249144 244682 249234
rect 244850 249144 245970 249234
rect 246138 249144 247902 249234
rect 248070 249144 248198 249234
rect 20 856 248198 249144
rect 130 734 1250 856
rect 1418 734 2538 856
rect 2706 734 4470 856
rect 4638 734 5758 856
rect 5926 734 7690 856
rect 7858 734 8978 856
rect 9146 734 10910 856
rect 11078 734 12198 856
rect 12366 734 14130 856
rect 14298 734 15418 856
rect 15586 734 17350 856
rect 17518 734 18638 856
rect 18806 734 20570 856
rect 20738 734 21858 856
rect 22026 734 23790 856
rect 23958 734 25078 856
rect 25246 734 27010 856
rect 27178 734 28298 856
rect 28466 734 30230 856
rect 30398 734 31518 856
rect 31686 734 33450 856
rect 33618 734 34738 856
rect 34906 734 36670 856
rect 36838 734 37958 856
rect 38126 734 39890 856
rect 40058 734 41178 856
rect 41346 734 43110 856
rect 43278 734 44398 856
rect 44566 734 46330 856
rect 46498 734 47618 856
rect 47786 734 49550 856
rect 49718 734 50838 856
rect 51006 734 52770 856
rect 52938 734 54058 856
rect 54226 734 55990 856
rect 56158 734 57278 856
rect 57446 734 59210 856
rect 59378 734 60498 856
rect 60666 734 62430 856
rect 62598 734 63718 856
rect 63886 734 65650 856
rect 65818 734 66938 856
rect 67106 734 68870 856
rect 69038 734 70158 856
rect 70326 734 72090 856
rect 72258 734 73378 856
rect 73546 734 75310 856
rect 75478 734 76598 856
rect 76766 734 78530 856
rect 78698 734 79818 856
rect 79986 734 81750 856
rect 81918 734 83038 856
rect 83206 734 84970 856
rect 85138 734 86258 856
rect 86426 734 88190 856
rect 88358 734 89478 856
rect 89646 734 91410 856
rect 91578 734 92698 856
rect 92866 734 94630 856
rect 94798 734 95918 856
rect 96086 734 97850 856
rect 98018 734 99138 856
rect 99306 734 101070 856
rect 101238 734 102358 856
rect 102526 734 104290 856
rect 104458 734 105578 856
rect 105746 734 107510 856
rect 107678 734 108798 856
rect 108966 734 110730 856
rect 110898 734 112018 856
rect 112186 734 113950 856
rect 114118 734 115238 856
rect 115406 734 117170 856
rect 117338 734 118458 856
rect 118626 734 120390 856
rect 120558 734 121678 856
rect 121846 734 123610 856
rect 123778 734 124898 856
rect 125066 734 126830 856
rect 126998 734 128118 856
rect 128286 734 130050 856
rect 130218 734 131338 856
rect 131506 734 133270 856
rect 133438 734 134558 856
rect 134726 734 136490 856
rect 136658 734 137778 856
rect 137946 734 139066 856
rect 139234 734 140998 856
rect 141166 734 142286 856
rect 142454 734 144218 856
rect 144386 734 145506 856
rect 145674 734 147438 856
rect 147606 734 148726 856
rect 148894 734 150658 856
rect 150826 734 151946 856
rect 152114 734 153878 856
rect 154046 734 155166 856
rect 155334 734 157098 856
rect 157266 734 158386 856
rect 158554 734 160318 856
rect 160486 734 161606 856
rect 161774 734 163538 856
rect 163706 734 164826 856
rect 164994 734 166758 856
rect 166926 734 168046 856
rect 168214 734 169978 856
rect 170146 734 171266 856
rect 171434 734 173198 856
rect 173366 734 174486 856
rect 174654 734 176418 856
rect 176586 734 177706 856
rect 177874 734 179638 856
rect 179806 734 180926 856
rect 181094 734 182858 856
rect 183026 734 184146 856
rect 184314 734 186078 856
rect 186246 734 187366 856
rect 187534 734 189298 856
rect 189466 734 190586 856
rect 190754 734 192518 856
rect 192686 734 193806 856
rect 193974 734 195738 856
rect 195906 734 197026 856
rect 197194 734 198958 856
rect 199126 734 200246 856
rect 200414 734 202178 856
rect 202346 734 203466 856
rect 203634 734 205398 856
rect 205566 734 206686 856
rect 206854 734 208618 856
rect 208786 734 209906 856
rect 210074 734 211838 856
rect 212006 734 213126 856
rect 213294 734 215058 856
rect 215226 734 216346 856
rect 216514 734 218278 856
rect 218446 734 219566 856
rect 219734 734 221498 856
rect 221666 734 222786 856
rect 222954 734 224718 856
rect 224886 734 226006 856
rect 226174 734 227938 856
rect 228106 734 229226 856
rect 229394 734 231158 856
rect 231326 734 232446 856
rect 232614 734 234378 856
rect 234546 734 235666 856
rect 235834 734 237598 856
rect 237766 734 238886 856
rect 239054 734 240818 856
rect 240986 734 242106 856
rect 242274 734 244038 856
rect 244206 734 245326 856
rect 245494 734 247258 856
rect 247426 734 248198 856
<< metal3 >>
rect 0 248888 800 249008
rect 249200 248888 250000 249008
rect 0 247528 800 247648
rect 249200 247528 250000 247648
rect 0 245488 800 245608
rect 249200 245488 250000 245608
rect 0 244128 800 244248
rect 249200 244128 250000 244248
rect 0 242088 800 242208
rect 249200 242088 250000 242208
rect 0 240728 800 240848
rect 249200 240728 250000 240848
rect 0 238688 800 238808
rect 249200 238688 250000 238808
rect 0 237328 800 237448
rect 249200 237328 250000 237448
rect 0 235288 800 235408
rect 249200 235288 250000 235408
rect 0 233928 800 234048
rect 249200 233928 250000 234048
rect 0 231888 800 232008
rect 249200 231888 250000 232008
rect 0 230528 800 230648
rect 249200 230528 250000 230648
rect 0 228488 800 228608
rect 249200 228488 250000 228608
rect 0 227128 800 227248
rect 249200 227128 250000 227248
rect 0 225088 800 225208
rect 249200 225088 250000 225208
rect 0 223728 800 223848
rect 249200 223728 250000 223848
rect 0 221688 800 221808
rect 249200 221688 250000 221808
rect 0 220328 800 220448
rect 249200 220328 250000 220448
rect 0 218288 800 218408
rect 249200 218288 250000 218408
rect 0 216928 800 217048
rect 249200 216928 250000 217048
rect 0 214888 800 215008
rect 249200 214888 250000 215008
rect 0 213528 800 213648
rect 249200 213528 250000 213648
rect 0 211488 800 211608
rect 249200 211488 250000 211608
rect 0 210128 800 210248
rect 249200 210128 250000 210248
rect 0 208088 800 208208
rect 249200 208088 250000 208208
rect 0 206728 800 206848
rect 249200 206728 250000 206848
rect 0 204688 800 204808
rect 249200 204688 250000 204808
rect 0 203328 800 203448
rect 249200 203328 250000 203448
rect 0 201288 800 201408
rect 249200 201288 250000 201408
rect 0 199928 800 200048
rect 249200 199928 250000 200048
rect 0 197888 800 198008
rect 249200 197888 250000 198008
rect 0 196528 800 196648
rect 249200 196528 250000 196648
rect 0 194488 800 194608
rect 249200 194488 250000 194608
rect 0 193128 800 193248
rect 249200 193128 250000 193248
rect 0 191088 800 191208
rect 249200 191088 250000 191208
rect 0 189728 800 189848
rect 249200 189728 250000 189848
rect 0 187688 800 187808
rect 249200 187688 250000 187808
rect 0 186328 800 186448
rect 249200 186328 250000 186448
rect 0 184288 800 184408
rect 249200 184288 250000 184408
rect 0 182928 800 183048
rect 249200 182928 250000 183048
rect 0 180888 800 181008
rect 249200 180888 250000 181008
rect 0 179528 800 179648
rect 249200 179528 250000 179648
rect 0 177488 800 177608
rect 249200 177488 250000 177608
rect 0 176128 800 176248
rect 249200 176128 250000 176248
rect 249200 174768 250000 174888
rect 0 174088 800 174208
rect 0 172728 800 172848
rect 249200 172728 250000 172848
rect 249200 171368 250000 171488
rect 0 170688 800 170808
rect 0 169328 800 169448
rect 249200 169328 250000 169448
rect 249200 167968 250000 168088
rect 0 167288 800 167408
rect 0 165928 800 166048
rect 249200 165928 250000 166048
rect 249200 164568 250000 164688
rect 0 163888 800 164008
rect 0 162528 800 162648
rect 249200 162528 250000 162648
rect 249200 161168 250000 161288
rect 0 160488 800 160608
rect 0 159128 800 159248
rect 249200 159128 250000 159248
rect 249200 157768 250000 157888
rect 0 157088 800 157208
rect 0 155728 800 155848
rect 249200 155728 250000 155848
rect 249200 154368 250000 154488
rect 0 153688 800 153808
rect 0 152328 800 152448
rect 249200 152328 250000 152448
rect 249200 150968 250000 151088
rect 0 150288 800 150408
rect 0 148928 800 149048
rect 249200 148928 250000 149048
rect 249200 147568 250000 147688
rect 0 146888 800 147008
rect 0 145528 800 145648
rect 249200 145528 250000 145648
rect 0 144168 800 144288
rect 249200 144168 250000 144288
rect 0 142128 800 142248
rect 249200 142128 250000 142248
rect 0 140768 800 140888
rect 249200 140768 250000 140888
rect 0 138728 800 138848
rect 249200 138728 250000 138848
rect 0 137368 800 137488
rect 249200 137368 250000 137488
rect 0 135328 800 135448
rect 249200 135328 250000 135448
rect 0 133968 800 134088
rect 249200 133968 250000 134088
rect 0 131928 800 132048
rect 249200 131928 250000 132048
rect 0 130568 800 130688
rect 249200 130568 250000 130688
rect 0 128528 800 128648
rect 249200 128528 250000 128648
rect 0 127168 800 127288
rect 249200 127168 250000 127288
rect 0 125128 800 125248
rect 249200 125128 250000 125248
rect 0 123768 800 123888
rect 249200 123768 250000 123888
rect 0 121728 800 121848
rect 249200 121728 250000 121848
rect 0 120368 800 120488
rect 249200 120368 250000 120488
rect 0 118328 800 118448
rect 249200 118328 250000 118448
rect 0 116968 800 117088
rect 249200 116968 250000 117088
rect 0 114928 800 115048
rect 249200 114928 250000 115048
rect 0 113568 800 113688
rect 249200 113568 250000 113688
rect 0 111528 800 111648
rect 249200 111528 250000 111648
rect 0 110168 800 110288
rect 249200 110168 250000 110288
rect 0 108128 800 108248
rect 249200 108128 250000 108248
rect 0 106768 800 106888
rect 249200 106768 250000 106888
rect 0 104728 800 104848
rect 249200 104728 250000 104848
rect 0 103368 800 103488
rect 249200 103368 250000 103488
rect 0 101328 800 101448
rect 249200 101328 250000 101448
rect 0 99968 800 100088
rect 249200 99968 250000 100088
rect 0 97928 800 98048
rect 249200 97928 250000 98048
rect 0 96568 800 96688
rect 249200 96568 250000 96688
rect 0 94528 800 94648
rect 249200 94528 250000 94648
rect 0 93168 800 93288
rect 249200 93168 250000 93288
rect 0 91128 800 91248
rect 249200 91128 250000 91248
rect 0 89768 800 89888
rect 249200 89768 250000 89888
rect 0 87728 800 87848
rect 249200 87728 250000 87848
rect 0 86368 800 86488
rect 249200 86368 250000 86488
rect 0 84328 800 84448
rect 249200 84328 250000 84448
rect 0 82968 800 83088
rect 249200 82968 250000 83088
rect 0 80928 800 81048
rect 249200 80928 250000 81048
rect 0 79568 800 79688
rect 249200 79568 250000 79688
rect 0 77528 800 77648
rect 249200 77528 250000 77648
rect 0 76168 800 76288
rect 249200 76168 250000 76288
rect 0 74128 800 74248
rect 249200 74128 250000 74248
rect 0 72768 800 72888
rect 249200 72768 250000 72888
rect 0 70728 800 70848
rect 249200 70728 250000 70848
rect 0 69368 800 69488
rect 249200 69368 250000 69488
rect 0 67328 800 67448
rect 249200 67328 250000 67448
rect 0 65968 800 66088
rect 249200 65968 250000 66088
rect 0 63928 800 64048
rect 249200 63928 250000 64048
rect 0 62568 800 62688
rect 249200 62568 250000 62688
rect 0 60528 800 60648
rect 249200 60528 250000 60648
rect 0 59168 800 59288
rect 249200 59168 250000 59288
rect 0 57128 800 57248
rect 249200 57128 250000 57248
rect 0 55768 800 55888
rect 249200 55768 250000 55888
rect 0 53728 800 53848
rect 249200 53728 250000 53848
rect 0 52368 800 52488
rect 249200 52368 250000 52488
rect 0 50328 800 50448
rect 249200 50328 250000 50448
rect 0 48968 800 49088
rect 249200 48968 250000 49088
rect 0 46928 800 47048
rect 249200 46928 250000 47048
rect 0 45568 800 45688
rect 249200 45568 250000 45688
rect 0 43528 800 43648
rect 249200 43528 250000 43648
rect 0 42168 800 42288
rect 249200 42168 250000 42288
rect 0 40128 800 40248
rect 249200 40128 250000 40248
rect 0 38768 800 38888
rect 249200 38768 250000 38888
rect 0 36728 800 36848
rect 249200 36728 250000 36848
rect 0 35368 800 35488
rect 249200 35368 250000 35488
rect 0 33328 800 33448
rect 249200 33328 250000 33448
rect 0 31968 800 32088
rect 249200 31968 250000 32088
rect 0 29928 800 30048
rect 249200 29928 250000 30048
rect 0 28568 800 28688
rect 249200 28568 250000 28688
rect 249200 27208 250000 27328
rect 0 26528 800 26648
rect 0 25168 800 25288
rect 249200 25168 250000 25288
rect 249200 23808 250000 23928
rect 0 23128 800 23248
rect 0 21768 800 21888
rect 249200 21768 250000 21888
rect 249200 20408 250000 20528
rect 0 19728 800 19848
rect 0 18368 800 18488
rect 249200 18368 250000 18488
rect 249200 17008 250000 17128
rect 0 16328 800 16448
rect 0 14968 800 15088
rect 249200 14968 250000 15088
rect 249200 13608 250000 13728
rect 0 12928 800 13048
rect 0 11568 800 11688
rect 249200 11568 250000 11688
rect 249200 10208 250000 10328
rect 0 9528 800 9648
rect 0 8168 800 8288
rect 249200 8168 250000 8288
rect 249200 6808 250000 6928
rect 0 6128 800 6248
rect 0 4768 800 4888
rect 249200 4768 250000 4888
rect 249200 3408 250000 3528
rect 0 2728 800 2848
rect 0 1368 800 1488
rect 249200 1368 250000 1488
rect 249200 8 250000 128
<< obsm3 >>
rect 880 248808 249120 248981
rect 800 247728 249200 248808
rect 880 247448 249120 247728
rect 800 245688 249200 247448
rect 880 245408 249120 245688
rect 800 244328 249200 245408
rect 880 244048 249120 244328
rect 800 242288 249200 244048
rect 880 242008 249120 242288
rect 800 240928 249200 242008
rect 880 240648 249120 240928
rect 800 238888 249200 240648
rect 880 238608 249120 238888
rect 800 237528 249200 238608
rect 880 237248 249120 237528
rect 800 235488 249200 237248
rect 880 235208 249120 235488
rect 800 234128 249200 235208
rect 880 233848 249120 234128
rect 800 232088 249200 233848
rect 880 231808 249120 232088
rect 800 230728 249200 231808
rect 880 230448 249120 230728
rect 800 228688 249200 230448
rect 880 228408 249120 228688
rect 800 227328 249200 228408
rect 880 227048 249120 227328
rect 800 225288 249200 227048
rect 880 225008 249120 225288
rect 800 223928 249200 225008
rect 880 223648 249120 223928
rect 800 221888 249200 223648
rect 880 221608 249120 221888
rect 800 220528 249200 221608
rect 880 220248 249120 220528
rect 800 218488 249200 220248
rect 880 218208 249120 218488
rect 800 217128 249200 218208
rect 880 216848 249120 217128
rect 800 215088 249200 216848
rect 880 214808 249120 215088
rect 800 213728 249200 214808
rect 880 213448 249120 213728
rect 800 211688 249200 213448
rect 880 211408 249120 211688
rect 800 210328 249200 211408
rect 880 210048 249120 210328
rect 800 208288 249200 210048
rect 880 208008 249120 208288
rect 800 206928 249200 208008
rect 880 206648 249120 206928
rect 800 204888 249200 206648
rect 880 204608 249120 204888
rect 800 203528 249200 204608
rect 880 203248 249120 203528
rect 800 201488 249200 203248
rect 880 201208 249120 201488
rect 800 200128 249200 201208
rect 880 199848 249120 200128
rect 800 198088 249200 199848
rect 880 197808 249120 198088
rect 800 196728 249200 197808
rect 880 196448 249120 196728
rect 800 194688 249200 196448
rect 880 194408 249120 194688
rect 800 193328 249200 194408
rect 880 193048 249120 193328
rect 800 191288 249200 193048
rect 880 191008 249120 191288
rect 800 189928 249200 191008
rect 880 189648 249120 189928
rect 800 187888 249200 189648
rect 880 187608 249120 187888
rect 800 186528 249200 187608
rect 880 186248 249120 186528
rect 800 184488 249200 186248
rect 880 184208 249120 184488
rect 800 183128 249200 184208
rect 880 182848 249120 183128
rect 800 181088 249200 182848
rect 880 180808 249120 181088
rect 800 179728 249200 180808
rect 880 179448 249120 179728
rect 800 177688 249200 179448
rect 880 177408 249120 177688
rect 800 176328 249200 177408
rect 880 176048 249120 176328
rect 800 174968 249200 176048
rect 800 174688 249120 174968
rect 800 174288 249200 174688
rect 880 174008 249200 174288
rect 800 172928 249200 174008
rect 880 172648 249120 172928
rect 800 171568 249200 172648
rect 800 171288 249120 171568
rect 800 170888 249200 171288
rect 880 170608 249200 170888
rect 800 169528 249200 170608
rect 880 169248 249120 169528
rect 800 168168 249200 169248
rect 800 167888 249120 168168
rect 800 167488 249200 167888
rect 880 167208 249200 167488
rect 800 166128 249200 167208
rect 880 165848 249120 166128
rect 800 164768 249200 165848
rect 800 164488 249120 164768
rect 800 164088 249200 164488
rect 880 163808 249200 164088
rect 800 162728 249200 163808
rect 880 162448 249120 162728
rect 800 161368 249200 162448
rect 800 161088 249120 161368
rect 800 160688 249200 161088
rect 880 160408 249200 160688
rect 800 159328 249200 160408
rect 880 159048 249120 159328
rect 800 157968 249200 159048
rect 800 157688 249120 157968
rect 800 157288 249200 157688
rect 880 157008 249200 157288
rect 800 155928 249200 157008
rect 880 155648 249120 155928
rect 800 154568 249200 155648
rect 800 154288 249120 154568
rect 800 153888 249200 154288
rect 880 153608 249200 153888
rect 800 152528 249200 153608
rect 880 152248 249120 152528
rect 800 151168 249200 152248
rect 800 150888 249120 151168
rect 800 150488 249200 150888
rect 880 150208 249200 150488
rect 800 149128 249200 150208
rect 880 148848 249120 149128
rect 800 147768 249200 148848
rect 800 147488 249120 147768
rect 800 147088 249200 147488
rect 880 146808 249200 147088
rect 800 145728 249200 146808
rect 880 145448 249120 145728
rect 800 144368 249200 145448
rect 880 144088 249120 144368
rect 800 142328 249200 144088
rect 880 142048 249120 142328
rect 800 140968 249200 142048
rect 880 140688 249120 140968
rect 800 138928 249200 140688
rect 880 138648 249120 138928
rect 800 137568 249200 138648
rect 880 137288 249120 137568
rect 800 135528 249200 137288
rect 880 135248 249120 135528
rect 800 134168 249200 135248
rect 880 133888 249120 134168
rect 800 132128 249200 133888
rect 880 131848 249120 132128
rect 800 130768 249200 131848
rect 880 130488 249120 130768
rect 800 128728 249200 130488
rect 880 128448 249120 128728
rect 800 127368 249200 128448
rect 880 127088 249120 127368
rect 800 125328 249200 127088
rect 880 125048 249120 125328
rect 800 123968 249200 125048
rect 880 123688 249120 123968
rect 800 121928 249200 123688
rect 880 121648 249120 121928
rect 800 120568 249200 121648
rect 880 120288 249120 120568
rect 800 118528 249200 120288
rect 880 118248 249120 118528
rect 800 117168 249200 118248
rect 880 116888 249120 117168
rect 800 115128 249200 116888
rect 880 114848 249120 115128
rect 800 113768 249200 114848
rect 880 113488 249120 113768
rect 800 111728 249200 113488
rect 880 111448 249120 111728
rect 800 110368 249200 111448
rect 880 110088 249120 110368
rect 800 108328 249200 110088
rect 880 108048 249120 108328
rect 800 106968 249200 108048
rect 880 106688 249120 106968
rect 800 104928 249200 106688
rect 880 104648 249120 104928
rect 800 103568 249200 104648
rect 880 103288 249120 103568
rect 800 101528 249200 103288
rect 880 101248 249120 101528
rect 800 100168 249200 101248
rect 880 99888 249120 100168
rect 800 98128 249200 99888
rect 880 97848 249120 98128
rect 800 96768 249200 97848
rect 880 96488 249120 96768
rect 800 94728 249200 96488
rect 880 94448 249120 94728
rect 800 93368 249200 94448
rect 880 93088 249120 93368
rect 800 91328 249200 93088
rect 880 91048 249120 91328
rect 800 89968 249200 91048
rect 880 89688 249120 89968
rect 800 87928 249200 89688
rect 880 87648 249120 87928
rect 800 86568 249200 87648
rect 880 86288 249120 86568
rect 800 84528 249200 86288
rect 880 84248 249120 84528
rect 800 83168 249200 84248
rect 880 82888 249120 83168
rect 800 81128 249200 82888
rect 880 80848 249120 81128
rect 800 79768 249200 80848
rect 880 79488 249120 79768
rect 800 77728 249200 79488
rect 880 77448 249120 77728
rect 800 76368 249200 77448
rect 880 76088 249120 76368
rect 800 74328 249200 76088
rect 880 74048 249120 74328
rect 800 72968 249200 74048
rect 880 72688 249120 72968
rect 800 70928 249200 72688
rect 880 70648 249120 70928
rect 800 69568 249200 70648
rect 880 69288 249120 69568
rect 800 67528 249200 69288
rect 880 67248 249120 67528
rect 800 66168 249200 67248
rect 880 65888 249120 66168
rect 800 64128 249200 65888
rect 880 63848 249120 64128
rect 800 62768 249200 63848
rect 880 62488 249120 62768
rect 800 60728 249200 62488
rect 880 60448 249120 60728
rect 800 59368 249200 60448
rect 880 59088 249120 59368
rect 800 57328 249200 59088
rect 880 57048 249120 57328
rect 800 55968 249200 57048
rect 880 55688 249120 55968
rect 800 53928 249200 55688
rect 880 53648 249120 53928
rect 800 52568 249200 53648
rect 880 52288 249120 52568
rect 800 50528 249200 52288
rect 880 50248 249120 50528
rect 800 49168 249200 50248
rect 880 48888 249120 49168
rect 800 47128 249200 48888
rect 880 46848 249120 47128
rect 800 45768 249200 46848
rect 880 45488 249120 45768
rect 800 43728 249200 45488
rect 880 43448 249120 43728
rect 800 42368 249200 43448
rect 880 42088 249120 42368
rect 800 40328 249200 42088
rect 880 40048 249120 40328
rect 800 38968 249200 40048
rect 880 38688 249120 38968
rect 800 36928 249200 38688
rect 880 36648 249120 36928
rect 800 35568 249200 36648
rect 880 35288 249120 35568
rect 800 33528 249200 35288
rect 880 33248 249120 33528
rect 800 32168 249200 33248
rect 880 31888 249120 32168
rect 800 30128 249200 31888
rect 880 29848 249120 30128
rect 800 28768 249200 29848
rect 880 28488 249120 28768
rect 800 27408 249200 28488
rect 800 27128 249120 27408
rect 800 26728 249200 27128
rect 880 26448 249200 26728
rect 800 25368 249200 26448
rect 880 25088 249120 25368
rect 800 24008 249200 25088
rect 800 23728 249120 24008
rect 800 23328 249200 23728
rect 880 23048 249200 23328
rect 800 21968 249200 23048
rect 880 21688 249120 21968
rect 800 20608 249200 21688
rect 800 20328 249120 20608
rect 800 19928 249200 20328
rect 880 19648 249200 19928
rect 800 18568 249200 19648
rect 880 18288 249120 18568
rect 800 17208 249200 18288
rect 800 16928 249120 17208
rect 800 16528 249200 16928
rect 880 16248 249200 16528
rect 800 15168 249200 16248
rect 880 14888 249120 15168
rect 800 13808 249200 14888
rect 800 13528 249120 13808
rect 800 13128 249200 13528
rect 880 12848 249200 13128
rect 800 11768 249200 12848
rect 880 11488 249120 11768
rect 800 10408 249200 11488
rect 800 10128 249120 10408
rect 800 9728 249200 10128
rect 880 9448 249200 9728
rect 800 8368 249200 9448
rect 880 8088 249120 8368
rect 800 7008 249200 8088
rect 800 6728 249120 7008
rect 800 6328 249200 6728
rect 880 6048 249200 6328
rect 800 4968 249200 6048
rect 880 4688 249120 4968
rect 800 3608 249200 4688
rect 800 3328 249120 3608
rect 800 2928 249200 3328
rect 880 2648 249200 2928
rect 800 1568 249200 2648
rect 880 1395 249120 1568
<< metal4 >>
rect 4208 2128 4528 247568
rect 19568 2128 19888 247568
rect 34928 2128 35248 247568
rect 50288 2128 50608 247568
rect 65648 2128 65968 247568
rect 81008 2128 81328 247568
rect 96368 2128 96688 247568
rect 111728 2128 112048 247568
rect 127088 2128 127408 247568
rect 142448 2128 142768 247568
rect 157808 2128 158128 247568
rect 173168 2128 173488 247568
rect 188528 2128 188848 247568
rect 203888 2128 204208 247568
rect 219248 2128 219568 247568
rect 234608 2128 234928 247568
<< obsm4 >>
rect 144683 97683 144749 99245
<< labels >>
rlabel metal2 s 238942 0 238998 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 249200 108128 250000 108248 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 85670 249200 85726 250000 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 249200 162528 250000 162648 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 72790 249200 72846 250000 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 249200 238688 250000 238808 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 93398 249200 93454 250000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 64418 249200 64474 250000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 77298 249200 77354 250000 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 249200 184288 250000 184408 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 11610 249200 11666 250000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 157798 249200 157854 250000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 69570 249200 69626 250000 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 114650 249200 114706 250000 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 0 210128 800 210248 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 170678 249200 170734 250000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 146850 249200 146906 250000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 249200 164568 250000 164688 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 236366 249200 236422 250000 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 249200 27208 250000 27328 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 249200 145528 250000 145648 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 121090 249200 121146 250000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 249200 86368 250000 86488 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 249200 80928 250000 81048 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 150070 249200 150126 250000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 88890 249200 88946 250000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 45098 249200 45154 250000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 249200 87728 250000 87848 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 3882 249200 3938 250000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 8390 249200 8446 250000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 164882 0 164938 800 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 47030 249200 47086 250000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 172610 249200 172666 250000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 249200 99968 250000 100088 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 249200 247528 250000 247648 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 199928 800 200048 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 30930 249200 30986 250000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 153290 249200 153346 250000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 249200 182928 250000 183048 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 249200 214888 250000 215008 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 225088 800 225208 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 34150 249200 34206 250000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 13542 249200 13598 250000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 48318 249200 48374 250000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 187688 800 187808 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 191286 249200 191342 250000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 180338 249200 180394 250000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 241518 249200 241574 250000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 27710 249200 27766 250000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 662 249200 718 250000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 235078 249200 235134 250000 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 249200 231888 250000 232008 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 249200 193128 250000 193248 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 249200 53728 250000 53848 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 249200 161168 250000 161288 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 249200 223728 250000 223848 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 249200 194488 250000 194608 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 247528 800 247648 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 232502 0 232558 800 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 249200 23808 250000 23928 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 174088 800 174208 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 51538 249200 51594 250000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 249200 137368 250000 137488 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 239586 249200 239642 250000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 249200 220328 250000 220448 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 249200 187688 250000 187808 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 247958 249200 248014 250000 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 249200 167968 250000 168088 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 50250 249200 50306 250000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 249200 20408 250000 20528 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 249200 154368 250000 154488 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 127530 249200 127586 250000 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 103058 249200 103114 250000 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 0 248888 800 249008 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 249200 97928 250000 98048 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 197726 249200 197782 250000 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 249200 125128 250000 125248 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 249200 67328 250000 67448 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 111430 249200 111486 250000 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 41878 249200 41934 250000 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 249200 228488 250000 228608 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 193128 800 193248 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 249200 155728 250000 155848 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 249200 21768 250000 21888 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 137190 249200 137246 250000 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 249200 62568 250000 62688 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 179050 249200 179106 250000 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 197888 800 198008 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 249200 157768 250000 157888 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 201288 800 201408 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 249200 35368 250000 35488 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 184846 249200 184902 250000 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 101770 249200 101826 250000 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 200946 249200 201002 250000 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 249200 148928 250000 149048 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 184288 800 184408 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 169390 249200 169446 250000 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 237654 0 237710 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 14830 249200 14886 250000 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 24490 249200 24546 250000 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 216402 0 216458 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 249200 179528 250000 179648 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 249200 103368 250000 103488 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 249200 210128 250000 210248 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 189998 249200 190054 250000 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 7102 249200 7158 250000 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 249200 130568 250000 130688 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 249200 45568 250000 45688 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 169328 800 169448 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 249200 199928 250000 200048 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 249200 147568 250000 147688 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 92110 249200 92166 250000 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 115938 249200 115994 250000 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 0 213528 800 213648 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 196438 249200 196494 250000 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 242806 249200 242862 250000 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 249200 106768 250000 106888 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 249200 111528 250000 111648 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 249200 191088 250000 191208 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 83738 249200 83794 250000 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 140768 800 140888 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 177118 249200 177174 250000 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 5170 249200 5226 250000 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 238298 249200 238354 250000 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 249200 43528 250000 43648 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 207386 249200 207442 250000 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 21270 249200 21326 250000 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 249200 57128 250000 57248 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 249200 235288 250000 235408 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 0 240728 800 240848 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 104990 249200 105046 250000 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 249200 180888 250000 181008 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 249200 96568 250000 96688 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 249200 59168 250000 59288 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 249200 42168 250000 42288 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 63130 249200 63186 250000 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 249200 159128 250000 159248 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 249200 197888 250000 198008 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 249200 65968 250000 66088 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 249200 74128 250000 74248 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 249200 76168 250000 76288 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 209318 249200 209374 250000 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 99838 249200 99894 250000 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 249200 176128 250000 176248 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 86958 249200 87014 250000 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 59910 249200 59966 250000 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 144918 249200 144974 250000 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 10322 249200 10378 250000 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 249200 8 250000 128 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 249200 17008 250000 17128 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 0 223728 800 223848 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 249200 114928 250000 115048 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 160488 800 160608 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 231858 249200 231914 250000 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 0 221688 800 221808 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 249200 89768 250000 89888 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 249200 133968 250000 134088 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 57978 249200 58034 250000 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 0 203328 800 203448 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 130750 249200 130806 250000 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 151358 249200 151414 250000 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 183558 249200 183614 250000 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 226706 249200 226762 250000 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 106278 249200 106334 250000 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 249200 218288 250000 218408 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 249200 52368 250000 52488 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 249200 3408 250000 3528 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 43810 249200 43866 250000 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 229926 249200 229982 250000 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 0 204688 800 204808 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 222842 0 222898 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 249200 221688 250000 221808 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 249200 110168 250000 110288 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 249200 121728 250000 121848 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 240874 0 240930 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 23202 249200 23258 250000 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 249200 38768 250000 38888 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 163888 800 164008 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 19982 249200 20038 250000 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 249200 242088 250000 242208 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 164238 249200 164294 250000 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 249200 91128 250000 91248 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 140410 249200 140466 250000 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 249200 113568 250000 113688 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 0 237328 800 237448 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 249200 31968 250000 32088 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 54758 249200 54814 250000 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 143630 249200 143686 250000 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 235722 0 235778 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 220266 249200 220322 250000 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 191088 800 191208 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 121728 800 121848 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 199658 249200 199714 250000 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 249200 63928 250000 64048 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 96618 249200 96674 250000 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 162528 800 162648 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 79230 249200 79286 250000 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 70858 249200 70914 250000 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 205454 0 205510 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 249200 1368 250000 1488 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 246026 249200 246082 250000 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 90178 249200 90234 250000 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 194488 800 194608 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 249200 123768 250000 123888 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 249200 116968 250000 117088 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 233146 249200 233202 250000 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 193218 249200 193274 250000 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 122378 249200 122434 250000 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 192574 0 192630 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 0 218288 800 218408 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 249200 131928 250000 132048 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 249200 50328 250000 50448 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 249200 28568 250000 28688 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 173254 0 173310 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 225418 249200 225474 250000 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 98550 249200 98606 250000 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 0 242088 800 242208 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 125598 249200 125654 250000 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 249200 18368 250000 18488 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 231214 0 231270 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 249200 48968 250000 49088 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 249200 36728 250000 36848 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 0 235288 800 235408 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 56690 249200 56746 250000 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 199014 0 199070 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 39302 249200 39358 250000 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 244094 0 244150 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 249200 127168 250000 127288 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 138478 249200 138534 250000 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 132038 249200 132094 250000 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 133970 249200 134026 250000 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 184202 0 184258 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 206742 0 206798 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 212538 249200 212594 250000 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 82450 249200 82506 250000 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 108210 249200 108266 250000 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 190642 0 190698 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 26422 249200 26478 250000 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 206098 249200 206154 250000 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 247314 0 247370 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 249200 245488 250000 245608 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 0 214888 800 215008 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 210606 249200 210662 250000 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 249200 142128 250000 142248 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 117870 249200 117926 250000 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 244738 249200 244794 250000 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 249200 138728 250000 138848 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 166170 249200 166226 250000 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 194506 249200 194562 250000 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 249200 189728 250000 189848 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 133968 800 134088 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 148138 249200 148194 250000 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 249200 237328 250000 237448 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 249200 94528 250000 94648 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 249200 140768 250000 140888 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 186328 800 186448 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 249200 206728 250000 206848 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 148928 800 149048 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 176128 800 176248 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 249200 60528 250000 60648 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 249200 171368 250000 171488 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 249200 40128 250000 40248 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 249200 33328 250000 33448 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 249200 233928 250000 234048 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 249200 101328 250000 101448 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 218978 249200 219034 250000 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 249200 135328 250000 135448 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 249246 249200 249302 250000 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 222198 249200 222254 250000 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 74078 249200 74134 250000 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 32862 249200 32918 250000 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 249200 77528 250000 77648 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 249200 144168 250000 144288 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 249200 203328 250000 203448 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 170688 800 170808 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 228638 249200 228694 250000 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 0 220328 800 220448 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 16762 249200 16818 250000 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 0 216928 800 217048 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 249200 11568 250000 11688 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 234434 0 234490 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 249200 72768 250000 72888 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 249200 204688 250000 204808 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 177488 800 177608 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 119158 249200 119214 250000 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 80518 249200 80574 250000 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 249200 230528 250000 230648 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 189728 800 189848 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 66350 249200 66406 250000 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 249200 201288 250000 201408 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 175830 249200 175886 250000 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 0 238688 800 238808 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 202878 249200 202934 250000 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 215758 249200 215814 250000 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 217046 249200 217102 250000 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 135258 249200 135314 250000 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 249200 46928 250000 47048 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 0 245488 800 245608 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 128818 249200 128874 250000 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 0 208088 800 208208 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 249200 172728 250000 172848 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 249200 227128 250000 227248 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 182928 800 183048 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 249200 25168 250000 25288 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 249200 213528 250000 213648 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 95330 249200 95386 250000 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 249200 177488 250000 177608 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 249200 55768 250000 55888 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 76010 249200 76066 250000 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 249200 4768 250000 4888 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 0 231888 800 232008 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 249200 211488 250000 211608 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 249200 8168 250000 8288 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 1950 249200 2006 250000 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 156510 249200 156566 250000 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 0 244128 800 244248 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 18050 249200 18106 250000 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 247568 6 vssd1
port 503 nsew ground input
rlabel metal3 s 249200 70728 250000 70848 6 wb_clk_i
port 504 nsew signal input
rlabel metal3 s 0 228488 800 228608 6 wb_rst_i
port 505 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 109498 249200 109554 250000 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 53470 249200 53526 250000 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal3 s 0 196528 800 196648 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal3 s 249200 225088 250000 225208 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal3 s 249200 208088 250000 208208 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal3 s 249200 104728 250000 104848 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal3 s 249200 6808 250000 6928 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 112718 249200 112774 250000 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 188066 249200 188122 250000 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 150714 0 150770 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 215114 0 215170 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal3 s 249200 79568 250000 79688 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal3 s 0 227128 800 227248 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 37370 249200 37426 250000 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal3 s 249200 174768 250000 174888 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 223486 249200 223542 250000 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 159730 249200 159786 250000 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal3 s 249200 128528 250000 128648 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 203522 0 203578 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 154578 249200 154634 250000 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 195794 0 195850 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal3 s 249200 10208 250000 10328 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal3 s 249200 84328 250000 84448 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 40590 249200 40646 250000 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal3 s 249200 248888 250000 249008 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal3 s 249200 150968 250000 151088 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 141698 249200 141754 250000 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 204166 249200 204222 250000 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal3 s 0 230528 800 230648 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal3 s 249200 169328 250000 169448 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 213826 249200 213882 250000 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal3 s 249200 216928 250000 217048 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal3 s 249200 93168 250000 93288 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 186778 249200 186834 250000 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 36082 249200 36138 250000 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal3 s 249200 165928 250000 166048 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal3 s 249200 82968 250000 83088 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal3 s 249200 13608 250000 13728 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal3 s 249200 118328 250000 118448 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 181626 249200 181682 250000 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal3 s 249200 240728 250000 240848 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal3 s 249200 14968 250000 15088 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal3 s 249200 152328 250000 152448 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal3 s 249200 244128 250000 244248 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 173898 249200 173954 250000 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal3 s 249200 29928 250000 30048 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 168102 0 168158 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal3 s 0 206728 800 206848 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 61198 249200 61254 250000 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 124310 249200 124366 250000 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 67638 249200 67694 250000 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 167458 249200 167514 250000 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal3 s 249200 69368 250000 69488 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal3 s 0 159128 800 159248 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal3 s 249200 196528 250000 196648 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal3 s 249200 186328 250000 186448 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 162950 249200 163006 250000 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 161018 249200 161074 250000 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal3 s 0 233928 800 234048 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 29642 249200 29698 250000 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 wbs_stb_i
port 608 nsew signal input
rlabel metal3 s 249200 120368 250000 120488 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 250000 250000
string LEFview TRUE
string GDS_FILE /home/shahid/caravel_user_project/openlane/user_proj_systollic/runs/user_proj_systollic/results/magic/user_proj_systollic.gds
string GDS_END 19016606
string GDS_START 523702
<< end >>

