magic
tech sky130A
magscale 1 2
timestamp 1667209117
<< locali >>
rect 200129 539903 200163 540005
rect 84025 538339 84059 539529
rect 185961 538475 185995 539801
rect 188537 539087 188571 539801
rect 201969 538815 202003 539937
rect 207213 538407 207247 539937
rect 218713 538407 218747 539937
rect 229753 539291 229787 539937
rect 245393 538951 245427 540005
rect 262229 539019 262263 540073
rect 268393 538611 268427 540005
rect 272901 538271 272935 540005
rect 287161 539223 287195 540005
rect 289829 539155 289863 540005
rect 300869 539019 300903 540073
rect 303445 538679 303479 540073
rect 320189 538679 320223 540073
rect 322765 538747 322799 540073
rect 328561 539155 328595 540073
rect 339509 538747 339543 540073
rect 355609 539359 355643 540073
rect 413569 538271 413603 540141
rect 416145 538543 416179 540141
rect 424517 538883 424551 540141
rect 57897 85459 57931 85969
rect 80069 60367 80103 60809
rect 143549 60435 143583 60877
rect 149161 60435 149195 60945
rect 168389 59891 168423 61285
rect 211077 59891 211111 61285
rect 218069 59891 218103 61217
rect 224693 59891 224727 61217
rect 236009 59823 236043 61013
rect 254041 59755 254075 61081
rect 257997 59755 258031 61081
rect 258089 59755 258123 61149
rect 286977 59755 287011 61149
rect 291117 59755 291151 61013
rect 302249 59755 302283 61761
rect 315957 59755 315991 61761
rect 350457 60503 350491 60945
rect 358829 59755 358863 61693
rect 375297 59687 375331 61693
rect 375389 59755 375423 61625
rect 378057 59755 378091 61625
rect 400137 59755 400171 60877
rect 404277 59755 404311 60809
rect 431877 59619 431911 60741
rect 125517 57715 125551 57749
rect 125517 57681 125793 57715
rect 139995 57681 140237 57715
rect 279525 57579 279559 57817
rect 409521 57239 409555 57613
rect 404461 56967 404495 57205
rect 388453 4471 388487 4981
rect 77309 3927 77343 4097
rect 100769 2975 100803 3621
rect 127633 3111 127667 3757
rect 307769 3383 307803 3825
rect 524337 3587 524371 3961
<< viali >>
rect 413569 540141 413603 540175
rect 262229 540073 262263 540107
rect 200129 540005 200163 540039
rect 245393 540005 245427 540039
rect 200129 539869 200163 539903
rect 201969 539937 202003 539971
rect 185961 539801 185995 539835
rect 84025 539529 84059 539563
rect 188537 539801 188571 539835
rect 188537 539053 188571 539087
rect 201969 538781 202003 538815
rect 207213 539937 207247 539971
rect 185961 538441 185995 538475
rect 207213 538373 207247 538407
rect 218713 539937 218747 539971
rect 229753 539937 229787 539971
rect 229753 539257 229787 539291
rect 300869 540073 300903 540107
rect 262229 538985 262263 539019
rect 268393 540005 268427 540039
rect 245393 538917 245427 538951
rect 268393 538577 268427 538611
rect 272901 540005 272935 540039
rect 218713 538373 218747 538407
rect 84025 538305 84059 538339
rect 287161 540005 287195 540039
rect 287161 539189 287195 539223
rect 289829 540005 289863 540039
rect 289829 539121 289863 539155
rect 300869 538985 300903 539019
rect 303445 540073 303479 540107
rect 303445 538645 303479 538679
rect 320189 540073 320223 540107
rect 322765 540073 322799 540107
rect 328561 540073 328595 540107
rect 328561 539121 328595 539155
rect 339509 540073 339543 540107
rect 322765 538713 322799 538747
rect 355609 540073 355643 540107
rect 355609 539325 355643 539359
rect 339509 538713 339543 538747
rect 320189 538645 320223 538679
rect 272901 538237 272935 538271
rect 416145 540141 416179 540175
rect 424517 540141 424551 540175
rect 424517 538849 424551 538883
rect 416145 538509 416179 538543
rect 413569 538237 413603 538271
rect 57897 85969 57931 86003
rect 57897 85425 57931 85459
rect 302249 61761 302283 61795
rect 168389 61285 168423 61319
rect 149161 60945 149195 60979
rect 143549 60877 143583 60911
rect 80069 60809 80103 60843
rect 143549 60401 143583 60435
rect 149161 60401 149195 60435
rect 80069 60333 80103 60367
rect 168389 59857 168423 59891
rect 211077 61285 211111 61319
rect 211077 59857 211111 59891
rect 218069 61217 218103 61251
rect 218069 59857 218103 59891
rect 224693 61217 224727 61251
rect 258089 61149 258123 61183
rect 254041 61081 254075 61115
rect 224693 59857 224727 59891
rect 236009 61013 236043 61047
rect 236009 59789 236043 59823
rect 254041 59721 254075 59755
rect 257997 61081 258031 61115
rect 257997 59721 258031 59755
rect 258089 59721 258123 59755
rect 286977 61149 287011 61183
rect 286977 59721 287011 59755
rect 291117 61013 291151 61047
rect 291117 59721 291151 59755
rect 302249 59721 302283 59755
rect 315957 61761 315991 61795
rect 358829 61693 358863 61727
rect 350457 60945 350491 60979
rect 350457 60469 350491 60503
rect 315957 59721 315991 59755
rect 358829 59721 358863 59755
rect 375297 61693 375331 61727
rect 375389 61625 375423 61659
rect 375389 59721 375423 59755
rect 378057 61625 378091 61659
rect 378057 59721 378091 59755
rect 400137 60877 400171 60911
rect 400137 59721 400171 59755
rect 404277 60809 404311 60843
rect 404277 59721 404311 59755
rect 431877 60741 431911 60775
rect 375297 59653 375331 59687
rect 431877 59585 431911 59619
rect 279525 57817 279559 57851
rect 125517 57749 125551 57783
rect 125793 57681 125827 57715
rect 139961 57681 139995 57715
rect 140237 57681 140271 57715
rect 279525 57545 279559 57579
rect 409521 57613 409555 57647
rect 404461 57205 404495 57239
rect 409521 57205 409555 57239
rect 404461 56933 404495 56967
rect 388453 4981 388487 5015
rect 388453 4437 388487 4471
rect 77309 4097 77343 4131
rect 77309 3893 77343 3927
rect 524337 3961 524371 3995
rect 307769 3825 307803 3859
rect 127633 3757 127667 3791
rect 100769 3621 100803 3655
rect 524337 3553 524371 3587
rect 307769 3349 307803 3383
rect 127633 3077 127667 3111
rect 100769 2941 100803 2975
<< metal1 >>
rect 144822 700816 144828 700868
rect 144880 700856 144886 700868
rect 170306 700856 170312 700868
rect 144880 700828 170312 700856
rect 144880 700816 144886 700828
rect 170306 700816 170312 700828
rect 170364 700816 170370 700868
rect 92382 700748 92388 700800
rect 92440 700788 92446 700800
rect 202782 700788 202788 700800
rect 92440 700760 202788 700788
rect 92440 700748 92446 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 57790 700680 57796 700732
rect 57848 700720 57854 700732
rect 154114 700720 154120 700732
rect 57848 700692 154120 700720
rect 57848 700680 57854 700692
rect 154114 700680 154120 700692
rect 154172 700680 154178 700732
rect 172422 700680 172428 700732
rect 172480 700720 172486 700732
rect 300118 700720 300124 700732
rect 172480 700692 300124 700720
rect 172480 700680 172486 700692
rect 300118 700680 300124 700692
rect 300176 700680 300182 700732
rect 122742 700612 122748 700664
rect 122800 700652 122806 700664
rect 235166 700652 235172 700664
rect 122800 700624 235172 700652
rect 122800 700612 122806 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 283834 700612 283840 700664
rect 283892 700652 283898 700664
rect 439498 700652 439504 700664
rect 283892 700624 439504 700652
rect 283892 700612 283898 700624
rect 439498 700612 439504 700624
rect 439556 700612 439562 700664
rect 137830 700544 137836 700596
rect 137888 700584 137894 700596
rect 304994 700584 305000 700596
rect 137888 700556 305000 700584
rect 137888 700544 137894 700556
rect 304994 700544 305000 700556
rect 305052 700544 305058 700596
rect 429838 700544 429844 700596
rect 429896 700584 429902 700596
rect 440418 700584 440424 700596
rect 429896 700556 440424 700584
rect 429896 700544 429902 700556
rect 440418 700544 440424 700556
rect 440476 700544 440482 700596
rect 57514 700476 57520 700528
rect 57572 700516 57578 700528
rect 332502 700516 332508 700528
rect 57572 700488 332508 700516
rect 57572 700476 57578 700488
rect 332502 700476 332508 700488
rect 332560 700476 332566 700528
rect 348786 700476 348792 700528
rect 348844 700516 348850 700528
rect 439866 700516 439872 700528
rect 348844 700488 439872 700516
rect 348844 700476 348850 700488
rect 439866 700476 439872 700488
rect 439924 700476 439930 700528
rect 464338 700476 464344 700528
rect 464396 700516 464402 700528
rect 478506 700516 478512 700528
rect 464396 700488 478512 700516
rect 464396 700476 464402 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 57606 700408 57612 700460
rect 57664 700448 57670 700460
rect 397454 700448 397460 700460
rect 57664 700420 397460 700448
rect 57664 700408 57670 700420
rect 397454 700408 397460 700420
rect 397512 700408 397518 700460
rect 413646 700408 413652 700460
rect 413704 700448 413710 700460
rect 439774 700448 439780 700460
rect 413704 700420 439780 700448
rect 413704 700408 413710 700420
rect 439774 700408 439780 700420
rect 439832 700408 439838 700460
rect 447778 700408 447784 700460
rect 447836 700448 447842 700460
rect 527174 700448 527180 700460
rect 447836 700420 527180 700448
rect 447836 700408 447842 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 59262 700340 59268 700392
rect 59320 700380 59326 700392
rect 72970 700380 72976 700392
rect 59320 700352 72976 700380
rect 59320 700340 59326 700352
rect 72970 700340 72976 700352
rect 73028 700340 73034 700392
rect 136542 700340 136548 700392
rect 136600 700380 136606 700392
rect 559650 700380 559656 700392
rect 136600 700352 559656 700380
rect 136600 700340 136606 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 440602 700312 440608 700324
rect 8168 700284 440608 700312
rect 8168 700272 8174 700284
rect 440602 700272 440608 700284
rect 440660 700272 440666 700324
rect 442350 700272 442356 700324
rect 442408 700312 442414 700324
rect 543458 700312 543464 700324
rect 442408 700284 543464 700312
rect 442408 700272 442414 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 48222 698912 48228 698964
rect 48280 698952 48286 698964
rect 494790 698952 494796 698964
rect 48280 698924 494796 698952
rect 48280 698912 48286 698924
rect 494790 698912 494796 698924
rect 494848 698912 494854 698964
rect 266354 697620 266360 697672
rect 266412 697660 266418 697672
rect 267642 697660 267648 697672
rect 266412 697632 267648 697660
rect 266412 697620 266418 697632
rect 267642 697620 267648 697632
rect 267700 697620 267706 697672
rect 89162 697552 89168 697604
rect 89220 697592 89226 697604
rect 449894 697592 449900 697604
rect 89220 697564 449900 697592
rect 89220 697552 89226 697564
rect 449894 697552 449900 697564
rect 449952 697552 449958 697604
rect 89622 696940 89628 696992
rect 89680 696980 89686 696992
rect 580166 696980 580172 696992
rect 89680 696952 580172 696980
rect 89680 696940 89686 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 440786 683176 440792 683188
rect 3476 683148 440792 683176
rect 3476 683136 3482 683148
rect 440786 683136 440792 683148
rect 440844 683136 440850 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 439406 670732 439412 670744
rect 3568 670704 439412 670732
rect 3568 670692 3574 670704
rect 439406 670692 439412 670704
rect 439464 670692 439470 670744
rect 442258 670692 442264 670744
rect 442316 670732 442322 670744
rect 580166 670732 580172 670744
rect 442316 670704 580172 670732
rect 442316 670692 442322 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 440326 656928 440332 656940
rect 3476 656900 440332 656928
rect 3476 656888 3482 656900
rect 440326 656888 440332 656900
rect 440384 656888 440390 656940
rect 57698 630640 57704 630692
rect 57756 630680 57762 630692
rect 580166 630680 580172 630692
rect 57756 630652 580172 630680
rect 57756 630640 57762 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 158622 616836 158628 616888
rect 158680 616876 158686 616888
rect 580166 616876 580172 616888
rect 158680 616848 580172 616876
rect 158680 616836 158686 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 164142 590656 164148 590708
rect 164200 590696 164206 590708
rect 579614 590696 579620 590708
rect 164200 590668 579620 590696
rect 164200 590656 164206 590668
rect 579614 590656 579620 590668
rect 579672 590656 579678 590708
rect 3510 579640 3516 579692
rect 3568 579680 3574 579692
rect 281534 579680 281540 579692
rect 3568 579652 281540 579680
rect 3568 579640 3574 579652
rect 281534 579640 281540 579652
rect 281592 579640 281598 579692
rect 442442 576852 442448 576904
rect 442500 576892 442506 576904
rect 579614 576892 579620 576904
rect 442500 576864 579620 576892
rect 442500 576852 442506 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 47946 563048 47952 563100
rect 48004 563088 48010 563100
rect 579890 563088 579896 563100
rect 48004 563060 579896 563088
rect 48004 563048 48010 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 91554 543532 91560 543584
rect 91612 543572 91618 543584
rect 92382 543572 92388 543584
rect 91612 543544 92388 543572
rect 91612 543532 91618 543544
rect 92382 543532 92388 543544
rect 92440 543532 92446 543584
rect 121822 543532 121828 543584
rect 121880 543572 121886 543584
rect 122742 543572 122748 543584
rect 121880 543544 122748 543572
rect 121880 543532 121886 543544
rect 122742 543532 122748 543544
rect 122800 543532 122806 543584
rect 157886 543532 157892 543584
rect 157944 543572 157950 543584
rect 158622 543572 158628 543584
rect 157944 543544 158628 543572
rect 157944 543532 157950 543544
rect 158622 543532 158628 543544
rect 158680 543532 158686 543584
rect 163038 543532 163044 543584
rect 163096 543572 163102 543584
rect 164142 543572 164148 543584
rect 163096 543544 164148 543572
rect 163096 543532 163102 543544
rect 164142 543532 164148 543544
rect 164200 543532 164206 543584
rect 171410 543532 171416 543584
rect 171468 543572 171474 543584
rect 172422 543572 172428 543584
rect 171468 543544 172428 543572
rect 171468 543532 171474 543544
rect 172422 543532 172428 543544
rect 172480 543532 172486 543584
rect 427078 543328 427084 543380
rect 427136 543368 427142 543380
rect 440510 543368 440516 543380
rect 427136 543340 440516 543368
rect 427136 543328 427142 543340
rect 440510 543328 440516 543340
rect 440568 543328 440574 543380
rect 4062 543260 4068 543312
rect 4120 543300 4126 543312
rect 80606 543300 80612 543312
rect 4120 543272 80612 543300
rect 4120 543260 4126 543272
rect 80606 543260 80612 543272
rect 80664 543260 80670 543312
rect 173986 543260 173992 543312
rect 174044 543300 174050 543312
rect 450078 543300 450084 543312
rect 174044 543272 450084 543300
rect 174044 543260 174050 543272
rect 450078 543260 450084 543272
rect 450136 543260 450142 543312
rect 29638 543192 29644 543244
rect 29696 543232 29702 543244
rect 94774 543232 94780 543244
rect 29696 543204 94780 543232
rect 29696 543192 29702 543204
rect 94774 543192 94780 543204
rect 94832 543192 94838 543244
rect 108298 543192 108304 543244
rect 108356 543232 108362 543244
rect 439590 543232 439596 543244
rect 108356 543204 439596 543232
rect 108356 543192 108362 543204
rect 439590 543192 439596 543204
rect 439648 543192 439654 543244
rect 16482 543124 16488 543176
rect 16540 543164 16546 543176
rect 61286 543164 61292 543176
rect 16540 543136 61292 543164
rect 16540 543124 16546 543136
rect 61286 543124 61292 543136
rect 61344 543124 61350 543176
rect 78030 543124 78036 543176
rect 78088 543164 78094 543176
rect 448606 543164 448612 543176
rect 78088 543136 448612 543164
rect 78088 543124 78094 543136
rect 448606 543124 448612 543136
rect 448664 543124 448670 543176
rect 3694 543056 3700 543108
rect 3752 543096 3758 543108
rect 64506 543096 64512 543108
rect 3752 543068 64512 543096
rect 3752 543056 3758 543068
rect 64506 543056 64512 543068
rect 64564 543056 64570 543108
rect 418706 543056 418712 543108
rect 418764 543096 418770 543108
rect 445846 543096 445852 543108
rect 418764 543068 445852 543096
rect 418764 543056 418770 543068
rect 445846 543056 445852 543068
rect 445904 543056 445910 543108
rect 3510 542988 3516 543040
rect 3568 543028 3574 543040
rect 99926 543028 99932 543040
rect 3568 543000 99932 543028
rect 3568 542988 3574 543000
rect 99926 542988 99932 543000
rect 99984 542988 99990 543040
rect 407758 542988 407764 543040
rect 407816 543028 407822 543040
rect 475378 543028 475384 543040
rect 407816 543000 475384 543028
rect 407816 542988 407822 543000
rect 475378 542988 475384 543000
rect 475436 542988 475442 543040
rect 48130 542920 48136 542972
rect 48188 542960 48194 542972
rect 102502 542960 102508 542972
rect 48188 542932 102508 542960
rect 48188 542920 48194 542932
rect 102502 542920 102508 542932
rect 102560 542920 102566 542972
rect 369762 542920 369768 542972
rect 369820 542960 369826 542972
rect 444374 542960 444380 542972
rect 369820 542932 444380 542960
rect 369820 542920 369826 542932
rect 444374 542920 444380 542932
rect 444432 542920 444438 542972
rect 8202 542852 8208 542904
rect 8260 542892 8266 542904
rect 199102 542892 199108 542904
rect 8260 542864 199108 542892
rect 8260 542852 8266 542864
rect 199102 542852 199108 542864
rect 199160 542852 199166 542904
rect 259638 542852 259644 542904
rect 259696 542892 259702 542904
rect 449986 542892 449992 542904
rect 259696 542864 449992 542892
rect 259696 542852 259702 542864
rect 449986 542852 449992 542864
rect 450044 542852 450050 542904
rect 12342 542784 12348 542836
rect 12400 542824 12406 542836
rect 204254 542824 204260 542836
rect 12400 542796 204260 542824
rect 12400 542784 12406 542796
rect 204254 542784 204260 542796
rect 204312 542784 204318 542836
rect 248690 542784 248696 542836
rect 248748 542824 248754 542836
rect 452654 542824 452660 542836
rect 248748 542796 452660 542824
rect 248748 542784 248754 542796
rect 452654 542784 452660 542796
rect 452712 542784 452718 542836
rect 27522 542716 27528 542768
rect 27580 542756 27586 542768
rect 275738 542756 275744 542768
rect 27580 542728 275744 542756
rect 27580 542716 27586 542728
rect 275738 542716 275744 542728
rect 275796 542716 275802 542768
rect 325326 542716 325332 542768
rect 325384 542756 325390 542768
rect 511258 542756 511264 542768
rect 325384 542728 511264 542756
rect 325384 542716 325390 542728
rect 511258 542716 511264 542728
rect 511316 542716 511322 542768
rect 25498 542648 25504 542700
rect 25556 542688 25562 542700
rect 97350 542688 97356 542700
rect 25556 542660 97356 542688
rect 25556 542648 25562 542660
rect 97350 542648 97356 542660
rect 97408 542648 97414 542700
rect 182358 542648 182364 542700
rect 182416 542688 182422 542700
rect 454126 542688 454132 542700
rect 182416 542660 454132 542688
rect 182416 542648 182422 542660
rect 454126 542648 454132 542660
rect 454184 542648 454190 542700
rect 56686 542580 56692 542632
rect 56744 542620 56750 542632
rect 333698 542620 333704 542632
rect 56744 542592 333704 542620
rect 56744 542580 56750 542592
rect 333698 542580 333704 542592
rect 333756 542580 333762 542632
rect 405182 542580 405188 542632
rect 405240 542620 405246 542632
rect 498838 542620 498844 542632
rect 405240 542592 498844 542620
rect 405240 542580 405246 542592
rect 498838 542580 498844 542592
rect 498896 542580 498902 542632
rect 3234 542512 3240 542564
rect 3292 542552 3298 542564
rect 130194 542552 130200 542564
rect 3292 542524 130200 542552
rect 3292 542512 3298 542524
rect 130194 542512 130200 542524
rect 130252 542512 130258 542564
rect 143718 542512 143724 542564
rect 143776 542552 143782 542564
rect 144822 542552 144828 542564
rect 143776 542524 144828 542552
rect 143776 542512 143782 542524
rect 144822 542512 144828 542524
rect 144880 542512 144886 542564
rect 55030 542444 55036 542496
rect 55088 542484 55094 542496
rect 67082 542484 67088 542496
rect 55088 542456 67088 542484
rect 55088 542444 55094 542456
rect 67082 542444 67088 542456
rect 67140 542444 67146 542496
rect 430298 542444 430304 542496
rect 430356 542484 430362 542496
rect 503714 542484 503720 542496
rect 430356 542456 503720 542484
rect 430356 542444 430362 542456
rect 503714 542444 503720 542456
rect 503772 542444 503778 542496
rect 54294 542376 54300 542428
rect 54352 542416 54358 542428
rect 69658 542416 69664 542428
rect 54352 542388 69664 542416
rect 54352 542376 54358 542388
rect 69658 542376 69664 542388
rect 69716 542376 69722 542428
rect 432874 542376 432880 542428
rect 432932 542416 432938 542428
rect 439682 542416 439688 542428
rect 432932 542388 439688 542416
rect 432932 542376 432938 542388
rect 439682 542376 439688 542388
rect 439740 542376 439746 542428
rect 45370 541628 45376 541680
rect 45428 541668 45434 541680
rect 266354 541668 266360 541680
rect 45428 541640 266360 541668
rect 45428 541628 45434 541640
rect 266354 541628 266360 541640
rect 266412 541628 266418 541680
rect 374914 541560 374920 541612
rect 374972 541600 374978 541612
rect 456978 541600 456984 541612
rect 374972 541572 456984 541600
rect 374972 541560 374978 541572
rect 456978 541560 456984 541572
rect 457036 541560 457042 541612
rect 372338 541492 372344 541544
rect 372396 541532 372402 541544
rect 479518 541532 479524 541544
rect 372396 541504 479524 541532
rect 372396 541492 372402 541504
rect 479518 541492 479524 541504
rect 479576 541492 479582 541544
rect 400030 541424 400036 541476
rect 400088 541464 400094 541476
rect 522298 541464 522304 541476
rect 400088 541436 522304 541464
rect 400088 541424 400094 541436
rect 522298 541424 522304 541436
rect 522356 541424 522362 541476
rect 344646 541356 344652 541408
rect 344704 541396 344710 541408
rect 486418 541396 486424 541408
rect 344704 541368 486424 541396
rect 344704 541356 344710 541368
rect 486418 541356 486424 541368
rect 486476 541356 486482 541408
rect 421926 541288 421932 541340
rect 421984 541328 421990 541340
rect 566458 541328 566464 541340
rect 421984 541300 566464 541328
rect 421984 541288 421990 541300
rect 566458 541288 566464 541300
rect 566516 541288 566522 541340
rect 237742 541220 237748 541272
rect 237800 541260 237806 541272
rect 454034 541260 454040 541272
rect 237800 541232 454040 541260
rect 237800 541220 237806 541232
rect 454034 541220 454040 541232
rect 454092 541220 454098 541272
rect 264790 541152 264796 541204
rect 264848 541192 264854 541204
rect 518158 541192 518164 541204
rect 264848 541164 518164 541192
rect 264848 541152 264854 541164
rect 518158 541152 518164 541164
rect 518216 541152 518222 541204
rect 196526 541084 196532 541136
rect 196584 541124 196590 541136
rect 458818 541124 458824 541136
rect 196584 541096 458824 541124
rect 196584 541084 196590 541096
rect 458818 541084 458824 541096
rect 458876 541084 458882 541136
rect 212626 541016 212632 541068
rect 212684 541056 212690 541068
rect 499574 541056 499580 541068
rect 212684 541028 499580 541056
rect 212684 541016 212690 541028
rect 499574 541016 499580 541028
rect 499632 541016 499638 541068
rect 152090 540948 152096 541000
rect 152148 540988 152154 541000
rect 456794 540988 456800 541000
rect 152148 540960 456800 540988
rect 152148 540948 152154 540960
rect 456794 540948 456800 540960
rect 456852 540948 456858 541000
rect 48038 540268 48044 540320
rect 48096 540308 48102 540320
rect 104894 540308 104900 540320
rect 48096 540280 104900 540308
rect 48096 540268 48102 540280
rect 104894 540268 104900 540280
rect 104952 540268 104958 540320
rect 49510 540200 49516 540252
rect 49568 540240 49574 540252
rect 364334 540240 364340 540252
rect 49568 540212 364340 540240
rect 49568 540200 49574 540212
rect 364334 540200 364340 540212
rect 364392 540200 364398 540252
rect 413554 540172 413560 540184
rect 413515 540144 413560 540172
rect 413554 540132 413560 540144
rect 413612 540132 413618 540184
rect 416130 540172 416136 540184
rect 416091 540144 416136 540172
rect 416130 540132 416136 540144
rect 416188 540132 416194 540184
rect 424502 540172 424508 540184
rect 424463 540144 424508 540172
rect 424502 540132 424508 540144
rect 424560 540132 424566 540184
rect 262214 540104 262220 540116
rect 262175 540076 262220 540104
rect 262214 540064 262220 540076
rect 262272 540064 262278 540116
rect 300854 540104 300860 540116
rect 300815 540076 300860 540104
rect 300854 540064 300860 540076
rect 300912 540064 300918 540116
rect 303430 540104 303436 540116
rect 303391 540076 303436 540104
rect 303430 540064 303436 540076
rect 303488 540064 303494 540116
rect 320174 540104 320180 540116
rect 320135 540076 320180 540104
rect 320174 540064 320180 540076
rect 320232 540064 320238 540116
rect 322750 540104 322756 540116
rect 322711 540076 322756 540104
rect 322750 540064 322756 540076
rect 322808 540064 322814 540116
rect 328546 540104 328552 540116
rect 328507 540076 328552 540104
rect 328546 540064 328552 540076
rect 328604 540064 328610 540116
rect 339494 540104 339500 540116
rect 339455 540076 339500 540104
rect 339494 540064 339500 540076
rect 339552 540064 339558 540116
rect 355594 540104 355600 540116
rect 355555 540076 355600 540104
rect 355594 540064 355600 540076
rect 355652 540064 355658 540116
rect 363966 540064 363972 540116
rect 364024 540104 364030 540116
rect 468478 540104 468484 540116
rect 364024 540076 468484 540104
rect 364024 540064 364030 540076
rect 468478 540064 468484 540076
rect 468536 540064 468542 540116
rect 200117 540039 200175 540045
rect 200117 540005 200129 540039
rect 200163 540036 200175 540039
rect 245378 540036 245384 540048
rect 200163 540008 209774 540036
rect 245339 540008 245384 540036
rect 200163 540005 200175 540008
rect 200117 539999 200175 540005
rect 193674 539928 193680 539980
rect 193732 539968 193738 539980
rect 201954 539968 201960 539980
rect 193732 539940 201724 539968
rect 201915 539940 201960 539968
rect 193732 539928 193738 539940
rect 141418 539860 141424 539912
rect 141476 539900 141482 539912
rect 200117 539903 200175 539909
rect 200117 539900 200129 539903
rect 141476 539872 200129 539900
rect 141476 539860 141482 539872
rect 200117 539869 200129 539872
rect 200163 539869 200175 539903
rect 200117 539863 200175 539869
rect 185946 539832 185952 539844
rect 185907 539804 185952 539832
rect 185946 539792 185952 539804
rect 186004 539792 186010 539844
rect 188522 539832 188528 539844
rect 188483 539804 188528 539832
rect 188522 539792 188528 539804
rect 188580 539792 188586 539844
rect 201696 539832 201724 539940
rect 201954 539928 201960 539940
rect 202012 539928 202018 539980
rect 207198 539968 207204 539980
rect 207159 539940 207204 539968
rect 207198 539928 207204 539940
rect 207256 539928 207262 539980
rect 209746 539900 209774 540008
rect 245378 539996 245384 540008
rect 245436 539996 245442 540048
rect 268378 540036 268384 540048
rect 268339 540008 268384 540036
rect 268378 539996 268384 540008
rect 268436 539996 268442 540048
rect 272886 540036 272892 540048
rect 272847 540008 272892 540036
rect 272886 539996 272892 540008
rect 272944 539996 272950 540048
rect 287146 540036 287152 540048
rect 287107 540008 287152 540036
rect 287146 539996 287152 540008
rect 287204 539996 287210 540048
rect 289814 540036 289820 540048
rect 289775 540008 289820 540036
rect 289814 539996 289820 540008
rect 289872 539996 289878 540048
rect 295242 539996 295248 540048
rect 295300 540036 295306 540048
rect 493318 540036 493324 540048
rect 295300 540008 493324 540036
rect 295300 539996 295306 540008
rect 493318 539996 493324 540008
rect 493376 539996 493382 540048
rect 218698 539968 218704 539980
rect 218659 539940 218704 539968
rect 218698 539928 218704 539940
rect 218756 539928 218762 539980
rect 229738 539968 229744 539980
rect 229699 539940 229744 539968
rect 229738 539928 229744 539940
rect 229796 539928 229802 539980
rect 234430 539928 234436 539980
rect 234488 539968 234494 539980
rect 513374 539968 513380 539980
rect 234488 539940 513380 539968
rect 234488 539928 234494 539940
rect 513374 539928 513380 539940
rect 513432 539928 513438 539980
rect 455414 539900 455420 539912
rect 209746 539872 455420 539900
rect 455414 539860 455420 539872
rect 455472 539860 455478 539912
rect 531406 539832 531412 539844
rect 201696 539804 531412 539832
rect 531406 539792 531412 539804
rect 531464 539792 531470 539844
rect 3326 539724 3332 539776
rect 3384 539764 3390 539776
rect 446030 539764 446036 539776
rect 3384 539736 446036 539764
rect 3384 539724 3390 539736
rect 446030 539724 446036 539736
rect 446088 539724 446094 539776
rect 111242 539656 111248 539708
rect 111300 539696 111306 539708
rect 502334 539696 502340 539708
rect 111300 539668 502340 539696
rect 111300 539656 111306 539668
rect 502334 539656 502340 539668
rect 502392 539656 502398 539708
rect 86770 539588 86776 539640
rect 86828 539628 86834 539640
rect 556246 539628 556252 539640
rect 86828 539600 556252 539628
rect 86828 539588 86834 539600
rect 556246 539588 556252 539600
rect 556304 539588 556310 539640
rect 84010 539560 84016 539572
rect 83971 539532 84016 539560
rect 84010 539520 84016 539532
rect 84068 539520 84074 539572
rect 160738 539520 160744 539572
rect 160796 539560 160802 539572
rect 160796 539532 437474 539560
rect 160796 539520 160802 539532
rect 4798 539452 4804 539504
rect 4856 539492 4862 539504
rect 435174 539492 435180 539504
rect 4856 539464 435180 539492
rect 4856 539452 4862 539464
rect 435174 539452 435180 539464
rect 435232 539452 435238 539504
rect 437446 539492 437474 539532
rect 438394 539520 438400 539572
rect 438452 539560 438458 539572
rect 442994 539560 443000 539572
rect 438452 539532 443000 539560
rect 438452 539520 438458 539532
rect 442994 539520 443000 539532
rect 443052 539520 443058 539572
rect 440234 539492 440240 539504
rect 437446 539464 440240 539492
rect 440234 539452 440240 539464
rect 440292 539452 440298 539504
rect 60642 539384 60648 539436
rect 60700 539424 60706 539436
rect 440970 539424 440976 539436
rect 60700 539396 440976 539424
rect 60700 539384 60706 539396
rect 440970 539384 440976 539396
rect 441028 539384 441034 539436
rect 355597 539359 355655 539365
rect 355597 539325 355609 539359
rect 355643 539356 355655 539359
rect 543734 539356 543740 539368
rect 355643 539328 543740 539356
rect 355643 539325 355655 539328
rect 355597 539319 355655 539325
rect 543734 539316 543740 539328
rect 543792 539316 543798 539368
rect 229741 539291 229799 539297
rect 229741 539257 229753 539291
rect 229787 539288 229799 539291
rect 441062 539288 441068 539300
rect 229787 539260 441068 539288
rect 229787 539257 229799 539260
rect 229741 539251 229799 539257
rect 441062 539248 441068 539260
rect 441120 539248 441126 539300
rect 46842 539180 46848 539232
rect 46900 539220 46906 539232
rect 287149 539223 287207 539229
rect 287149 539220 287161 539223
rect 46900 539192 287161 539220
rect 46900 539180 46906 539192
rect 287149 539189 287161 539192
rect 287195 539189 287207 539223
rect 287149 539183 287207 539189
rect 316954 539180 316960 539232
rect 317012 539220 317018 539232
rect 511994 539220 512000 539232
rect 317012 539192 512000 539220
rect 317012 539180 317018 539192
rect 511994 539180 512000 539192
rect 512052 539180 512058 539232
rect 44082 539112 44088 539164
rect 44140 539152 44146 539164
rect 289817 539155 289875 539161
rect 289817 539152 289829 539155
rect 44140 539124 289829 539152
rect 44140 539112 44146 539124
rect 289817 539121 289829 539124
rect 289863 539121 289875 539155
rect 289817 539115 289875 539121
rect 328549 539155 328607 539161
rect 328549 539121 328561 539155
rect 328595 539152 328607 539155
rect 529934 539152 529940 539164
rect 328595 539124 529940 539152
rect 328595 539121 328607 539124
rect 328549 539115 328607 539121
rect 529934 539112 529940 539124
rect 529992 539112 529998 539164
rect 188525 539087 188583 539093
rect 188525 539053 188537 539087
rect 188571 539084 188583 539087
rect 440878 539084 440884 539096
rect 188571 539056 440884 539084
rect 188571 539053 188583 539056
rect 188525 539047 188583 539053
rect 440878 539044 440884 539056
rect 440936 539044 440942 539096
rect 3510 538976 3516 539028
rect 3568 539016 3574 539028
rect 262217 539019 262275 539025
rect 262217 539016 262229 539019
rect 3568 538988 262229 539016
rect 3568 538976 3574 538988
rect 262217 538985 262229 538988
rect 262263 538985 262275 539019
rect 262217 538979 262275 538985
rect 300857 539019 300915 539025
rect 300857 538985 300869 539019
rect 300903 539016 300915 539019
rect 550634 539016 550640 539028
rect 300903 538988 550640 539016
rect 300903 538985 300915 538988
rect 300857 538979 300915 538985
rect 550634 538976 550640 538988
rect 550692 538976 550698 539028
rect 245381 538951 245439 538957
rect 245381 538917 245393 538951
rect 245427 538948 245439 538951
rect 505094 538948 505100 538960
rect 245427 538920 505100 538948
rect 245427 538917 245439 538920
rect 245381 538911 245439 538917
rect 505094 538908 505100 538920
rect 505152 538908 505158 538960
rect 424505 538883 424563 538889
rect 424505 538849 424517 538883
rect 424551 538880 424563 538883
rect 580166 538880 580172 538892
rect 424551 538852 580172 538880
rect 424551 538849 424563 538852
rect 424505 538843 424563 538849
rect 580166 538840 580172 538852
rect 580224 538840 580230 538892
rect 201957 538815 202015 538821
rect 201957 538781 201969 538815
rect 202003 538812 202015 538815
rect 483014 538812 483020 538824
rect 202003 538784 483020 538812
rect 202003 538781 202015 538784
rect 201957 538775 202015 538781
rect 483014 538772 483020 538784
rect 483072 538772 483078 538824
rect 38562 538704 38568 538756
rect 38620 538744 38626 538756
rect 322753 538747 322811 538753
rect 322753 538744 322765 538747
rect 38620 538716 322765 538744
rect 38620 538704 38626 538716
rect 322753 538713 322765 538716
rect 322799 538713 322811 538747
rect 322753 538707 322811 538713
rect 339497 538747 339555 538753
rect 339497 538713 339509 538747
rect 339543 538744 339555 538747
rect 580534 538744 580540 538756
rect 339543 538716 580540 538744
rect 339543 538713 339555 538716
rect 339497 538707 339555 538713
rect 580534 538704 580540 538716
rect 580592 538704 580598 538756
rect 3878 538636 3884 538688
rect 3936 538676 3942 538688
rect 303433 538679 303491 538685
rect 303433 538676 303445 538679
rect 3936 538648 303445 538676
rect 3936 538636 3942 538648
rect 303433 538645 303445 538648
rect 303479 538645 303491 538679
rect 303433 538639 303491 538645
rect 320177 538679 320235 538685
rect 320177 538645 320189 538679
rect 320223 538676 320235 538679
rect 580902 538676 580908 538688
rect 320223 538648 580908 538676
rect 320223 538645 320235 538648
rect 320177 538639 320235 538645
rect 580902 538636 580908 538648
rect 580960 538636 580966 538688
rect 268381 538611 268439 538617
rect 268381 538577 268393 538611
rect 268427 538608 268439 538611
rect 580718 538608 580724 538620
rect 268427 538580 580724 538608
rect 268427 538577 268439 538580
rect 268381 538571 268439 538577
rect 580718 538568 580724 538580
rect 580776 538568 580782 538620
rect 416133 538543 416191 538549
rect 416133 538509 416145 538543
rect 416179 538540 416191 538543
rect 580626 538540 580632 538552
rect 416179 538512 580632 538540
rect 416179 538509 416191 538512
rect 416133 538503 416191 538509
rect 580626 538500 580632 538512
rect 580684 538500 580690 538552
rect 185949 538475 186007 538481
rect 185949 538441 185961 538475
rect 185995 538472 186007 538475
rect 539686 538472 539692 538484
rect 185995 538444 539692 538472
rect 185995 538441 186007 538444
rect 185949 538435 186007 538441
rect 539686 538432 539692 538444
rect 539744 538432 539750 538484
rect 3694 538364 3700 538416
rect 3752 538404 3758 538416
rect 207201 538407 207259 538413
rect 207201 538404 207213 538407
rect 3752 538376 207213 538404
rect 3752 538364 3758 538376
rect 207201 538373 207213 538376
rect 207247 538373 207259 538407
rect 207201 538367 207259 538373
rect 218701 538407 218759 538413
rect 218701 538373 218713 538407
rect 218747 538404 218759 538407
rect 580074 538404 580080 538416
rect 218747 538376 580080 538404
rect 218747 538373 218759 538376
rect 218701 538367 218759 538373
rect 580074 538364 580080 538376
rect 580132 538364 580138 538416
rect 84013 538339 84071 538345
rect 84013 538305 84025 538339
rect 84059 538336 84071 538339
rect 487154 538336 487160 538348
rect 84059 538308 487160 538336
rect 84059 538305 84071 538308
rect 84013 538299 84071 538305
rect 487154 538296 487160 538308
rect 487212 538296 487218 538348
rect 3970 538228 3976 538280
rect 4028 538268 4034 538280
rect 272889 538271 272947 538277
rect 272889 538268 272901 538271
rect 4028 538240 272901 538268
rect 4028 538228 4034 538240
rect 272889 538237 272901 538240
rect 272935 538237 272947 538271
rect 272889 538231 272947 538237
rect 413557 538271 413615 538277
rect 413557 538237 413569 538271
rect 413603 538268 413615 538271
rect 580442 538268 580448 538280
rect 413603 538240 580448 538268
rect 413603 538237 413615 538240
rect 413557 538231 413615 538237
rect 580442 538228 580448 538240
rect 580500 538228 580506 538280
rect 59814 537888 59820 537940
rect 59872 537928 59878 537940
rect 466454 537928 466460 537940
rect 59872 537900 466460 537928
rect 59872 537888 59878 537900
rect 466454 537888 466460 537900
rect 466512 537888 466518 537940
rect 9582 537820 9588 537872
rect 9640 537860 9646 537872
rect 439958 537860 439964 537872
rect 9640 537832 439964 537860
rect 9640 537820 9646 537832
rect 439958 537820 439964 537832
rect 440016 537820 440022 537872
rect 57330 537752 57336 537804
rect 57388 537792 57394 537804
rect 580902 537792 580908 537804
rect 57388 537764 580908 537792
rect 57388 537752 57394 537764
rect 580902 537752 580908 537764
rect 580960 537752 580966 537804
rect 442074 531292 442080 531344
rect 442132 531332 442138 531344
rect 481634 531332 481640 531344
rect 442132 531304 481640 531332
rect 442132 531292 442138 531304
rect 481634 531292 481640 531304
rect 481692 531292 481698 531344
rect 55122 529932 55128 529984
rect 55180 529972 55186 529984
rect 57422 529972 57428 529984
rect 55180 529944 57428 529972
rect 55180 529932 55186 529944
rect 57422 529932 57428 529944
rect 57480 529932 57486 529984
rect 43990 527144 43996 527196
rect 44048 527184 44054 527196
rect 57330 527184 57336 527196
rect 44048 527156 57336 527184
rect 44048 527144 44054 527156
rect 57330 527144 57336 527156
rect 57388 527144 57394 527196
rect 54938 524424 54944 524476
rect 54996 524464 55002 524476
rect 57330 524464 57336 524476
rect 54996 524436 57336 524464
rect 54996 524424 55002 524436
rect 57330 524424 57336 524436
rect 57388 524424 57394 524476
rect 442534 523608 442540 523660
rect 442592 523648 442598 523660
rect 448514 523648 448520 523660
rect 442592 523620 448520 523648
rect 442592 523608 442598 523620
rect 448514 523608 448520 523620
rect 448572 523608 448578 523660
rect 50982 520276 50988 520328
rect 51040 520316 51046 520328
rect 57330 520316 57336 520328
rect 51040 520288 57336 520316
rect 51040 520276 51046 520288
rect 57330 520276 57336 520288
rect 57388 520276 57394 520328
rect 52362 517488 52368 517540
rect 52420 517528 52426 517540
rect 57330 517528 57336 517540
rect 52420 517500 57336 517528
rect 52420 517488 52426 517500
rect 57330 517488 57336 517500
rect 57388 517488 57394 517540
rect 442902 517488 442908 517540
rect 442960 517528 442966 517540
rect 527818 517528 527824 517540
rect 442960 517500 527824 517528
rect 442960 517488 442966 517500
rect 527818 517488 527824 517500
rect 527876 517488 527882 517540
rect 46750 514768 46756 514820
rect 46808 514808 46814 514820
rect 57330 514808 57336 514820
rect 46808 514780 57336 514808
rect 46808 514768 46814 514780
rect 57330 514768 57336 514780
rect 57388 514768 57394 514820
rect 442902 514768 442908 514820
rect 442960 514808 442966 514820
rect 451274 514808 451280 514820
rect 442960 514780 451280 514808
rect 442960 514768 442966 514780
rect 451274 514768 451280 514780
rect 451332 514768 451338 514820
rect 442902 512184 442908 512236
rect 442960 512224 442966 512236
rect 445938 512224 445944 512236
rect 442960 512196 445944 512224
rect 442960 512184 442966 512196
rect 445938 512184 445944 512196
rect 445996 512184 446002 512236
rect 18598 511980 18604 512032
rect 18656 512020 18662 512032
rect 57330 512020 57336 512032
rect 18656 511992 57336 512020
rect 18656 511980 18662 511992
rect 57330 511980 57336 511992
rect 57388 511980 57394 512032
rect 3418 510552 3424 510604
rect 3476 510592 3482 510604
rect 57146 510592 57152 510604
rect 3476 510564 57152 510592
rect 3476 510552 3482 510564
rect 57146 510552 57152 510564
rect 57204 510552 57210 510604
rect 442534 505112 442540 505164
rect 442592 505152 442598 505164
rect 447134 505152 447140 505164
rect 442592 505124 447140 505152
rect 442592 505112 442598 505124
rect 447134 505112 447140 505124
rect 447192 505112 447198 505164
rect 442810 502324 442816 502376
rect 442868 502364 442874 502376
rect 490006 502364 490012 502376
rect 442868 502336 490012 502364
rect 442868 502324 442874 502336
rect 490006 502324 490012 502336
rect 490064 502324 490070 502376
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 17218 501004 17224 501016
rect 3384 500976 17224 501004
rect 3384 500964 3390 500976
rect 17218 500964 17224 500976
rect 17276 500964 17282 501016
rect 442534 496816 442540 496868
rect 442592 496856 442598 496868
rect 447502 496856 447508 496868
rect 442592 496828 447508 496856
rect 442592 496816 442598 496828
rect 447502 496816 447508 496828
rect 447560 496816 447566 496868
rect 50890 491308 50896 491360
rect 50948 491348 50954 491360
rect 57606 491348 57612 491360
rect 50948 491320 57612 491348
rect 50948 491308 50954 491320
rect 57606 491308 57612 491320
rect 57664 491308 57670 491360
rect 45462 488520 45468 488572
rect 45520 488560 45526 488572
rect 57606 488560 57612 488572
rect 45520 488532 57612 488560
rect 45520 488520 45526 488532
rect 57606 488520 57612 488532
rect 57664 488520 57670 488572
rect 442718 485800 442724 485852
rect 442776 485840 442782 485852
rect 533338 485840 533344 485852
rect 442776 485812 533344 485840
rect 442776 485800 442782 485812
rect 533338 485800 533344 485812
rect 533396 485800 533402 485852
rect 52086 480224 52092 480276
rect 52144 480264 52150 480276
rect 57606 480264 57612 480276
rect 52144 480236 57612 480264
rect 52144 480224 52150 480236
rect 57606 480224 57612 480236
rect 57664 480224 57670 480276
rect 442902 480224 442908 480276
rect 442960 480264 442966 480276
rect 454678 480264 454684 480276
rect 442960 480236 454684 480264
rect 442960 480224 442966 480236
rect 454678 480224 454684 480236
rect 454736 480224 454742 480276
rect 50798 477504 50804 477556
rect 50856 477544 50862 477556
rect 57054 477544 57060 477556
rect 50856 477516 57060 477544
rect 50856 477504 50862 477516
rect 57054 477504 57060 477516
rect 57112 477504 57118 477556
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 14458 474756 14464 474768
rect 3476 474728 14464 474756
rect 3476 474716 3482 474728
rect 14458 474716 14464 474728
rect 14516 474716 14522 474768
rect 53742 474716 53748 474768
rect 53800 474756 53806 474768
rect 57606 474756 57612 474768
rect 53800 474728 57612 474756
rect 53800 474716 53806 474728
rect 57606 474716 57612 474728
rect 57664 474716 57670 474768
rect 442902 473356 442908 473408
rect 442960 473396 442966 473408
rect 456886 473396 456892 473408
rect 442960 473368 456892 473396
rect 442960 473356 442966 473368
rect 456886 473356 456892 473368
rect 456944 473356 456950 473408
rect 442902 470568 442908 470620
rect 442960 470608 442966 470620
rect 452746 470608 452752 470620
rect 442960 470580 452752 470608
rect 442960 470568 442966 470580
rect 452746 470568 452752 470580
rect 452804 470568 452810 470620
rect 51994 469208 52000 469260
rect 52052 469248 52058 469260
rect 57606 469248 57612 469260
rect 52052 469220 57612 469248
rect 52052 469208 52058 469220
rect 57606 469208 57612 469220
rect 57664 469208 57670 469260
rect 442902 468664 442908 468716
rect 442960 468704 442966 468716
rect 447594 468704 447600 468716
rect 442960 468676 447600 468704
rect 442960 468664 442966 468676
rect 447594 468664 447600 468676
rect 447652 468664 447658 468716
rect 54846 465060 54852 465112
rect 54904 465100 54910 465112
rect 56870 465100 56876 465112
rect 54904 465072 56876 465100
rect 54904 465060 54910 465072
rect 56870 465060 56876 465072
rect 56928 465060 56934 465112
rect 442810 465060 442816 465112
rect 442868 465100 442874 465112
rect 538858 465100 538864 465112
rect 442868 465072 538864 465100
rect 442868 465060 442874 465072
rect 538858 465060 538864 465072
rect 538916 465060 538922 465112
rect 442902 462544 442908 462596
rect 442960 462584 442966 462596
rect 447226 462584 447232 462596
rect 442960 462556 447232 462584
rect 442960 462544 442966 462556
rect 447226 462544 447232 462556
rect 447284 462544 447290 462596
rect 53650 462340 53656 462392
rect 53708 462380 53714 462392
rect 57606 462380 57612 462392
rect 53708 462352 57612 462380
rect 53708 462340 53714 462352
rect 57606 462340 57612 462352
rect 57664 462340 57670 462392
rect 442902 459824 442908 459876
rect 442960 459864 442966 459876
rect 447410 459864 447416 459876
rect 442960 459836 447416 459864
rect 442960 459824 442966 459836
rect 447410 459824 447416 459836
rect 447468 459824 447474 459876
rect 12250 459552 12256 459604
rect 12308 459592 12314 459604
rect 57606 459592 57612 459604
rect 12308 459564 57612 459592
rect 12308 459552 12314 459564
rect 57606 459552 57612 459564
rect 57664 459552 57670 459604
rect 442902 457104 442908 457156
rect 442960 457144 442966 457156
rect 447318 457144 447324 457156
rect 442960 457116 447324 457144
rect 442960 457104 442966 457116
rect 447318 457104 447324 457116
rect 447376 457104 447382 457156
rect 50706 456764 50712 456816
rect 50764 456804 50770 456816
rect 57606 456804 57612 456816
rect 50764 456776 57612 456804
rect 50764 456764 50770 456776
rect 57606 456764 57612 456776
rect 57664 456764 57670 456816
rect 54662 454044 54668 454096
rect 54720 454084 54726 454096
rect 57606 454084 57612 454096
rect 54720 454056 57612 454084
rect 54720 454044 54726 454056
rect 57606 454044 57612 454056
rect 57664 454044 57670 454096
rect 442902 454044 442908 454096
rect 442960 454084 442966 454096
rect 452838 454084 452844 454096
rect 442960 454056 452844 454084
rect 442960 454044 442966 454056
rect 452838 454044 452844 454056
rect 452896 454044 452902 454096
rect 2682 451256 2688 451308
rect 2740 451296 2746 451308
rect 57606 451296 57612 451308
rect 2740 451268 57612 451296
rect 2740 451256 2746 451268
rect 57606 451256 57612 451268
rect 57664 451256 57670 451308
rect 442902 447448 442908 447500
rect 442960 447488 442966 447500
rect 448698 447488 448704 447500
rect 442960 447460 448704 447488
rect 442960 447448 442966 447460
rect 448698 447448 448704 447460
rect 448756 447448 448762 447500
rect 3970 444388 3976 444440
rect 4028 444428 4034 444440
rect 57054 444428 57060 444440
rect 4028 444400 57060 444428
rect 4028 444388 4034 444400
rect 57054 444388 57060 444400
rect 57112 444388 57118 444440
rect 52270 436092 52276 436144
rect 52328 436132 52334 436144
rect 57606 436132 57612 436144
rect 52328 436104 57612 436132
rect 52328 436092 52334 436104
rect 57606 436092 57612 436104
rect 57664 436092 57670 436144
rect 442718 436092 442724 436144
rect 442776 436132 442782 436144
rect 516778 436132 516784 436144
rect 442776 436104 516784 436132
rect 442776 436092 442782 436104
rect 516778 436092 516784 436104
rect 516836 436092 516842 436144
rect 53558 433304 53564 433356
rect 53616 433344 53622 433356
rect 57606 433344 57612 433356
rect 53616 433316 57612 433344
rect 53616 433304 53622 433316
rect 57606 433304 57612 433316
rect 57664 433304 57670 433356
rect 440970 431876 440976 431928
rect 441028 431916 441034 431928
rect 579982 431916 579988 431928
rect 441028 431888 579988 431916
rect 441028 431876 441034 431888
rect 579982 431876 579988 431888
rect 580040 431876 580046 431928
rect 52178 430584 52184 430636
rect 52236 430624 52242 430636
rect 57606 430624 57612 430636
rect 52236 430596 57612 430624
rect 52236 430584 52242 430596
rect 57606 430584 57612 430596
rect 57664 430584 57670 430636
rect 442902 430584 442908 430636
rect 442960 430624 442966 430636
rect 448790 430624 448796 430636
rect 442960 430596 448796 430624
rect 442960 430584 442966 430596
rect 448790 430584 448796 430596
rect 448848 430584 448854 430636
rect 53374 427796 53380 427848
rect 53432 427836 53438 427848
rect 57606 427836 57612 427848
rect 53432 427808 57612 427836
rect 53432 427796 53438 427808
rect 57606 427796 57612 427808
rect 57664 427796 57670 427848
rect 5442 422288 5448 422340
rect 5500 422328 5506 422340
rect 57606 422328 57612 422340
rect 5500 422300 57612 422328
rect 5500 422288 5506 422300
rect 57606 422288 57612 422300
rect 57664 422288 57670 422340
rect 442902 422288 442908 422340
rect 442960 422328 442966 422340
rect 452930 422328 452936 422340
rect 442960 422300 452936 422328
rect 442960 422288 442966 422300
rect 452930 422288 452936 422300
rect 452988 422288 452994 422340
rect 46658 419500 46664 419552
rect 46716 419540 46722 419552
rect 57606 419540 57612 419552
rect 46716 419512 57612 419540
rect 46716 419500 46722 419512
rect 57606 419500 57612 419512
rect 57664 419500 57670 419552
rect 442534 418888 442540 418940
rect 442592 418928 442598 418940
rect 450170 418928 450176 418940
rect 442592 418900 450176 418928
rect 442592 418888 442598 418900
rect 450170 418888 450176 418900
rect 450228 418888 450234 418940
rect 50614 416780 50620 416832
rect 50672 416820 50678 416832
rect 57606 416820 57612 416832
rect 50672 416792 57612 416820
rect 50672 416780 50678 416792
rect 57606 416780 57612 416792
rect 57664 416780 57670 416832
rect 442718 415624 442724 415676
rect 442776 415664 442782 415676
rect 447686 415664 447692 415676
rect 442776 415636 447692 415664
rect 442776 415624 442782 415636
rect 447686 415624 447692 415636
rect 447744 415624 447750 415676
rect 54754 409844 54760 409896
rect 54812 409884 54818 409896
rect 57514 409884 57520 409896
rect 54812 409856 57520 409884
rect 54812 409844 54818 409856
rect 57514 409844 57520 409856
rect 57572 409844 57578 409896
rect 442534 409844 442540 409896
rect 442592 409884 442598 409896
rect 457070 409884 457076 409896
rect 442592 409856 457076 409884
rect 442592 409844 442598 409856
rect 457070 409844 457076 409856
rect 457128 409844 457134 409896
rect 442534 404608 442540 404660
rect 442592 404648 442598 404660
rect 446122 404648 446128 404660
rect 442592 404620 446128 404648
rect 442592 404608 442598 404620
rect 446122 404608 446128 404620
rect 446180 404608 446186 404660
rect 3602 402908 3608 402960
rect 3660 402948 3666 402960
rect 57514 402948 57520 402960
rect 3660 402920 57520 402948
rect 3660 402908 3666 402920
rect 57514 402908 57520 402920
rect 57572 402908 57578 402960
rect 49602 398828 49608 398880
rect 49660 398868 49666 398880
rect 57514 398868 57520 398880
rect 49660 398840 57520 398868
rect 49660 398828 49666 398840
rect 57514 398828 57520 398840
rect 57572 398828 57578 398880
rect 54202 396040 54208 396092
rect 54260 396080 54266 396092
rect 57514 396080 57520 396092
rect 54260 396052 57520 396080
rect 54260 396040 54266 396052
rect 57514 396040 57520 396052
rect 57572 396040 57578 396092
rect 442902 394952 442908 395004
rect 442960 394992 442966 395004
rect 448882 394992 448888 395004
rect 442960 394964 448888 394992
rect 442960 394952 442966 394964
rect 448882 394952 448888 394964
rect 448940 394952 448946 395004
rect 53466 393320 53472 393372
rect 53524 393360 53530 393372
rect 57514 393360 57520 393372
rect 53524 393332 57520 393360
rect 53524 393320 53530 393332
rect 57514 393320 57520 393332
rect 57572 393320 57578 393372
rect 47854 389172 47860 389224
rect 47912 389212 47918 389224
rect 57514 389212 57520 389224
rect 47912 389184 57520 389212
rect 47912 389172 47918 389184
rect 57514 389172 57520 389184
rect 57572 389172 57578 389224
rect 54478 387812 54484 387864
rect 54536 387852 54542 387864
rect 57514 387852 57520 387864
rect 54536 387824 57520 387852
rect 54536 387812 54542 387824
rect 57514 387812 57520 387824
rect 57572 387812 57578 387864
rect 51902 385024 51908 385076
rect 51960 385064 51966 385076
rect 57514 385064 57520 385076
rect 51960 385036 57520 385064
rect 51960 385024 51966 385036
rect 57514 385024 57520 385036
rect 57572 385024 57578 385076
rect 39298 380876 39304 380928
rect 39356 380916 39362 380928
rect 57514 380916 57520 380928
rect 39356 380888 57520 380916
rect 39356 380876 39362 380888
rect 57514 380876 57520 380888
rect 57572 380876 57578 380928
rect 442902 380876 442908 380928
rect 442960 380916 442966 380928
rect 518894 380916 518900 380928
rect 442960 380888 518900 380916
rect 442960 380876 442966 380888
rect 518894 380876 518900 380888
rect 518952 380876 518958 380928
rect 53098 378156 53104 378208
rect 53156 378196 53162 378208
rect 57514 378196 57520 378208
rect 53156 378168 57520 378196
rect 53156 378156 53162 378168
rect 57514 378156 57520 378168
rect 57572 378156 57578 378208
rect 442902 378156 442908 378208
rect 442960 378196 442966 378208
rect 498194 378196 498200 378208
rect 442960 378168 498200 378196
rect 442960 378156 442966 378168
rect 498194 378156 498200 378168
rect 498252 378156 498258 378208
rect 442902 375368 442908 375420
rect 442960 375408 442966 375420
rect 508498 375408 508504 375420
rect 442960 375380 508504 375408
rect 442960 375368 442966 375380
rect 508498 375368 508504 375380
rect 508556 375368 508562 375420
rect 442902 372784 442908 372836
rect 442960 372824 442966 372836
rect 448974 372824 448980 372836
rect 442960 372796 448980 372824
rect 442960 372784 442966 372796
rect 448974 372784 448980 372796
rect 449032 372784 449038 372836
rect 50522 372580 50528 372632
rect 50580 372620 50586 372632
rect 57514 372620 57520 372632
rect 50580 372592 57520 372620
rect 50580 372580 50586 372592
rect 57514 372580 57520 372592
rect 57572 372580 57578 372632
rect 51534 367072 51540 367124
rect 51592 367112 51598 367124
rect 56870 367112 56876 367124
rect 51592 367084 56876 367112
rect 51592 367072 51598 367084
rect 56870 367072 56876 367084
rect 56928 367072 56934 367124
rect 442902 365712 442908 365764
rect 442960 365752 442966 365764
rect 547874 365752 547880 365764
rect 442960 365724 547880 365752
rect 442960 365712 442966 365724
rect 547874 365712 547880 365724
rect 547932 365712 547938 365764
rect 440878 365644 440884 365696
rect 440936 365684 440942 365696
rect 579982 365684 579988 365696
rect 440936 365656 579988 365684
rect 440936 365644 440942 365656
rect 579982 365644 579988 365656
rect 580040 365644 580046 365696
rect 51810 364352 51816 364404
rect 51868 364392 51874 364404
rect 56870 364392 56876 364404
rect 51868 364364 56876 364392
rect 51868 364352 51874 364364
rect 56870 364352 56876 364364
rect 56928 364352 56934 364404
rect 51718 361564 51724 361616
rect 51776 361604 51782 361616
rect 57514 361604 57520 361616
rect 51776 361576 57520 361604
rect 51776 361564 51782 361576
rect 57514 361564 57520 361576
rect 57572 361564 57578 361616
rect 442626 360544 442632 360596
rect 442684 360584 442690 360596
rect 443638 360584 443644 360596
rect 442684 360556 443644 360584
rect 442684 360544 442690 360556
rect 443638 360544 443644 360556
rect 443696 360544 443702 360596
rect 3786 358708 3792 358760
rect 3844 358748 3850 358760
rect 57514 358748 57520 358760
rect 3844 358720 57520 358748
rect 3844 358708 3850 358720
rect 57514 358708 57520 358720
rect 57572 358708 57578 358760
rect 442718 358368 442724 358420
rect 442776 358408 442782 358420
rect 447870 358408 447876 358420
rect 442776 358380 447876 358408
rect 442776 358368 442782 358380
rect 447870 358368 447876 358380
rect 447928 358368 447934 358420
rect 442902 354696 442908 354748
rect 442960 354736 442966 354748
rect 496814 354736 496820 354748
rect 442960 354708 496820 354736
rect 442960 354696 442966 354708
rect 496814 354696 496820 354708
rect 496872 354696 496878 354748
rect 442902 352384 442908 352436
rect 442960 352424 442966 352436
rect 444558 352424 444564 352436
rect 442960 352396 444564 352424
rect 442960 352384 442966 352396
rect 444558 352384 444564 352396
rect 444616 352384 444622 352436
rect 51626 351908 51632 351960
rect 51684 351948 51690 351960
rect 57514 351948 57520 351960
rect 51684 351920 57520 351948
rect 51684 351908 51690 351920
rect 57514 351908 57520 351920
rect 57572 351908 57578 351960
rect 45278 349120 45284 349172
rect 45336 349160 45342 349172
rect 56870 349160 56876 349172
rect 45336 349132 56876 349160
rect 45336 349120 45342 349132
rect 56870 349120 56876 349132
rect 56928 349120 56934 349172
rect 442718 349120 442724 349172
rect 442776 349160 442782 349172
rect 506566 349160 506572 349172
rect 442776 349132 506572 349160
rect 442776 349120 442782 349132
rect 506566 349120 506572 349132
rect 506624 349120 506630 349172
rect 54018 346400 54024 346452
rect 54076 346440 54082 346452
rect 57514 346440 57520 346452
rect 54076 346412 57520 346440
rect 54076 346400 54082 346412
rect 57514 346400 57520 346412
rect 57572 346400 57578 346452
rect 442902 342592 442908 342644
rect 442960 342632 442966 342644
rect 446306 342632 446312 342644
rect 442960 342604 446312 342632
rect 442960 342592 442966 342604
rect 446306 342592 446312 342604
rect 446364 342592 446370 342644
rect 54570 340892 54576 340944
rect 54628 340932 54634 340944
rect 57514 340932 57520 340944
rect 54628 340904 57520 340932
rect 54628 340892 54634 340904
rect 57514 340892 57520 340904
rect 57572 340892 57578 340944
rect 442902 340892 442908 340944
rect 442960 340932 442966 340944
rect 461578 340932 461584 340944
rect 442960 340904 461584 340932
rect 442960 340892 442966 340904
rect 461578 340892 461584 340904
rect 461636 340892 461642 340944
rect 53282 338104 53288 338156
rect 53340 338144 53346 338156
rect 57514 338144 57520 338156
rect 53340 338116 57520 338144
rect 53340 338104 53346 338116
rect 57514 338104 57520 338116
rect 57572 338104 57578 338156
rect 442902 338104 442908 338156
rect 442960 338144 442966 338156
rect 444650 338144 444656 338156
rect 442960 338116 444656 338144
rect 442960 338104 442966 338116
rect 444650 338104 444656 338116
rect 444708 338104 444714 338156
rect 442718 334160 442724 334212
rect 442776 334200 442782 334212
rect 446214 334200 446220 334212
rect 442776 334172 446220 334200
rect 442776 334160 442782 334172
rect 446214 334160 446220 334172
rect 446272 334160 446278 334212
rect 442902 331576 442908 331628
rect 442960 331616 442966 331628
rect 447962 331616 447968 331628
rect 442960 331588 447968 331616
rect 442960 331576 442966 331588
rect 447962 331576 447968 331588
rect 448020 331576 448026 331628
rect 53190 329808 53196 329860
rect 53248 329848 53254 329860
rect 57514 329848 57520 329860
rect 53248 329820 57520 329848
rect 53248 329808 53254 329820
rect 57514 329808 57520 329820
rect 57572 329808 57578 329860
rect 57514 329196 57520 329248
rect 57572 329236 57578 329248
rect 57882 329236 57888 329248
rect 57572 329208 57888 329236
rect 57572 329196 57578 329208
rect 57882 329196 57888 329208
rect 57940 329196 57946 329248
rect 442902 328448 442908 328500
rect 442960 328488 442966 328500
rect 454218 328488 454224 328500
rect 442960 328460 454224 328488
rect 442960 328448 442966 328460
rect 454218 328448 454224 328460
rect 454276 328448 454282 328500
rect 442534 326068 442540 326120
rect 442592 326108 442598 326120
rect 450262 326108 450268 326120
rect 442592 326080 450268 326108
rect 442592 326068 442598 326080
rect 450262 326068 450268 326080
rect 450320 326068 450326 326120
rect 442534 323076 442540 323128
rect 442592 323116 442598 323128
rect 443546 323116 443552 323128
rect 442592 323088 443552 323116
rect 442592 323076 442598 323088
rect 443546 323076 443552 323088
rect 443604 323076 443610 323128
rect 54386 322940 54392 322992
rect 54444 322980 54450 322992
rect 57330 322980 57336 322992
rect 54444 322952 57336 322980
rect 54444 322940 54450 322952
rect 57330 322940 57336 322952
rect 57388 322940 57394 322992
rect 442902 320152 442908 320204
rect 442960 320192 442966 320204
rect 451366 320192 451372 320204
rect 442960 320164 451372 320192
rect 442960 320152 442966 320164
rect 451366 320152 451372 320164
rect 451424 320152 451430 320204
rect 442902 317500 442908 317552
rect 442960 317540 442966 317552
rect 449066 317540 449072 317552
rect 442960 317512 449072 317540
rect 442960 317500 442966 317512
rect 449066 317500 449072 317512
rect 449124 317500 449130 317552
rect 52822 314644 52828 314696
rect 52880 314684 52886 314696
rect 56870 314684 56876 314696
rect 52880 314656 56876 314684
rect 52880 314644 52886 314656
rect 56870 314644 56876 314656
rect 56928 314644 56934 314696
rect 49418 311856 49424 311908
rect 49476 311896 49482 311908
rect 57330 311896 57336 311908
rect 49476 311868 57336 311896
rect 49476 311856 49482 311868
rect 57330 311856 57336 311868
rect 57388 311856 57394 311908
rect 442718 310768 442724 310820
rect 442776 310808 442782 310820
rect 444466 310808 444472 310820
rect 442776 310780 444472 310808
rect 442776 310768 442782 310780
rect 444466 310768 444472 310780
rect 444524 310768 444530 310820
rect 53006 309136 53012 309188
rect 53064 309176 53070 309188
rect 57330 309176 57336 309188
rect 53064 309148 57336 309176
rect 53064 309136 53070 309148
rect 57330 309136 57336 309148
rect 57388 309136 57394 309188
rect 442902 307776 442908 307828
rect 442960 307816 442966 307828
rect 465718 307816 465724 307828
rect 442960 307788 465724 307816
rect 442960 307776 442966 307788
rect 465718 307776 465724 307788
rect 465776 307776 465782 307828
rect 442442 302472 442448 302524
rect 442500 302512 442506 302524
rect 443270 302512 443276 302524
rect 442500 302484 443276 302512
rect 442500 302472 442506 302484
rect 443270 302472 443276 302484
rect 443328 302472 443334 302524
rect 43898 299480 43904 299532
rect 43956 299520 43962 299532
rect 57330 299520 57336 299532
rect 43956 299492 57336 299520
rect 43956 299480 43962 299492
rect 57330 299480 57336 299492
rect 57388 299480 57394 299532
rect 442902 298052 442908 298104
rect 442960 298092 442966 298104
rect 580902 298092 580908 298104
rect 442960 298064 580908 298092
rect 442960 298052 442966 298064
rect 580902 298052 580908 298064
rect 580960 298052 580966 298104
rect 21358 296692 21364 296744
rect 21416 296732 21422 296744
rect 57330 296732 57336 296744
rect 21416 296704 57336 296732
rect 21416 296692 21422 296704
rect 57330 296692 57336 296704
rect 57388 296692 57394 296744
rect 442442 294584 442448 294636
rect 442500 294624 442506 294636
rect 443362 294624 443368 294636
rect 442500 294596 443368 294624
rect 442500 294584 442506 294596
rect 443362 294584 443368 294596
rect 443420 294584 443426 294636
rect 47762 293972 47768 294024
rect 47820 294012 47826 294024
rect 57882 294012 57888 294024
rect 47820 293984 57888 294012
rect 47820 293972 47826 293984
rect 57882 293972 57888 293984
rect 57940 293972 57946 294024
rect 51258 291184 51264 291236
rect 51316 291224 51322 291236
rect 57054 291224 57060 291236
rect 51316 291196 57060 291224
rect 51316 291184 51322 291196
rect 57054 291184 57060 291196
rect 57112 291184 57118 291236
rect 442902 291184 442908 291236
rect 442960 291224 442966 291236
rect 448054 291224 448060 291236
rect 442960 291196 448060 291224
rect 442960 291184 442966 291196
rect 448054 291184 448060 291196
rect 448112 291184 448118 291236
rect 442902 288464 442908 288516
rect 442960 288504 442966 288516
rect 450354 288504 450360 288516
rect 442960 288476 450360 288504
rect 442960 288464 442966 288476
rect 450354 288464 450360 288476
rect 450412 288464 450418 288516
rect 52730 288396 52736 288448
rect 52788 288436 52794 288448
rect 57330 288436 57336 288448
rect 52788 288408 57336 288436
rect 52788 288396 52794 288408
rect 57330 288396 57336 288408
rect 57388 288396 57394 288448
rect 442902 285744 442908 285796
rect 442960 285784 442966 285796
rect 446398 285784 446404 285796
rect 442960 285756 446404 285784
rect 442960 285744 442966 285756
rect 446398 285744 446404 285756
rect 446456 285744 446462 285796
rect 50430 282888 50436 282940
rect 50488 282928 50494 282940
rect 57330 282928 57336 282940
rect 50488 282900 57336 282928
rect 50488 282888 50494 282900
rect 57330 282888 57336 282900
rect 57388 282888 57394 282940
rect 442810 278740 442816 278792
rect 442868 278780 442874 278792
rect 520918 278780 520924 278792
rect 442868 278752 520924 278780
rect 442868 278740 442874 278752
rect 520918 278740 520924 278752
rect 520976 278740 520982 278792
rect 51442 277380 51448 277432
rect 51500 277420 51506 277432
rect 57330 277420 57336 277432
rect 51500 277392 57336 277420
rect 51500 277380 51506 277392
rect 57330 277380 57336 277392
rect 57388 277380 57394 277432
rect 442534 276632 442540 276684
rect 442592 276672 442598 276684
rect 443454 276672 443460 276684
rect 442592 276644 443460 276672
rect 442592 276632 442598 276644
rect 443454 276632 443460 276644
rect 443512 276632 443518 276684
rect 442902 273232 442908 273284
rect 442960 273272 442966 273284
rect 529198 273272 529204 273284
rect 442960 273244 529204 273272
rect 442960 273232 442966 273244
rect 529198 273232 529204 273244
rect 529256 273232 529262 273284
rect 442902 270784 442908 270836
rect 442960 270824 442966 270836
rect 448238 270824 448244 270836
rect 442960 270796 448244 270824
rect 442960 270784 442966 270796
rect 448238 270784 448244 270796
rect 448296 270784 448302 270836
rect 52638 270512 52644 270564
rect 52696 270552 52702 270564
rect 57330 270552 57336 270564
rect 52696 270524 57336 270552
rect 52696 270512 52702 270524
rect 57330 270512 57336 270524
rect 57388 270512 57394 270564
rect 55674 268064 55680 268116
rect 55732 268104 55738 268116
rect 56594 268104 56600 268116
rect 55732 268076 56600 268104
rect 55732 268064 55738 268076
rect 56594 268064 56600 268076
rect 56652 268064 56658 268116
rect 442902 267724 442908 267776
rect 442960 267764 442966 267776
rect 454310 267764 454316 267776
rect 442960 267736 454316 267764
rect 442960 267724 442966 267736
rect 454310 267724 454316 267736
rect 454368 267724 454374 267776
rect 52914 264936 52920 264988
rect 52972 264976 52978 264988
rect 57422 264976 57428 264988
rect 52972 264948 57428 264976
rect 52972 264936 52978 264948
rect 57422 264936 57428 264948
rect 57480 264936 57486 264988
rect 442902 264936 442908 264988
rect 442960 264976 442966 264988
rect 485038 264976 485044 264988
rect 442960 264948 485044 264976
rect 442960 264936 442966 264948
rect 485038 264936 485044 264948
rect 485096 264936 485102 264988
rect 442902 263168 442908 263220
rect 442960 263208 442966 263220
rect 447778 263208 447784 263220
rect 442960 263180 447784 263208
rect 442960 263168 442966 263180
rect 447778 263168 447784 263180
rect 447836 263168 447842 263220
rect 51350 262216 51356 262268
rect 51408 262256 51414 262268
rect 57422 262256 57428 262268
rect 51408 262228 57428 262256
rect 51408 262216 51414 262228
rect 57422 262216 57428 262228
rect 57480 262216 57486 262268
rect 441062 259360 441068 259412
rect 441120 259400 441126 259412
rect 579798 259400 579804 259412
rect 441120 259372 579804 259400
rect 441120 259360 441126 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 442902 258068 442908 258120
rect 442960 258108 442966 258120
rect 472618 258108 472624 258120
rect 442960 258080 472624 258108
rect 442960 258068 442966 258080
rect 472618 258068 472624 258080
rect 472676 258068 472682 258120
rect 442534 256504 442540 256556
rect 442592 256544 442598 256556
rect 448146 256544 448152 256556
rect 442592 256516 448152 256544
rect 442592 256504 442598 256516
rect 448146 256504 448152 256516
rect 448204 256504 448210 256556
rect 2774 254056 2780 254108
rect 2832 254096 2838 254108
rect 4890 254096 4896 254108
rect 2832 254068 4896 254096
rect 2832 254056 2838 254068
rect 4890 254056 4896 254068
rect 4948 254056 4954 254108
rect 45186 253920 45192 253972
rect 45244 253960 45250 253972
rect 57422 253960 57428 253972
rect 45244 253932 57428 253960
rect 45244 253920 45250 253932
rect 57422 253920 57428 253932
rect 57480 253920 57486 253972
rect 442902 251132 442908 251184
rect 442960 251172 442966 251184
rect 580810 251172 580816 251184
rect 442960 251144 580816 251172
rect 442960 251132 442966 251144
rect 580810 251132 580816 251144
rect 580868 251132 580874 251184
rect 43806 249772 43812 249824
rect 43864 249812 43870 249824
rect 56870 249812 56876 249824
rect 43864 249784 56876 249812
rect 43864 249772 43870 249784
rect 56870 249772 56876 249784
rect 56928 249772 56934 249824
rect 442718 247052 442724 247104
rect 442776 247092 442782 247104
rect 454402 247092 454408 247104
rect 442776 247064 454408 247092
rect 442776 247052 442782 247064
rect 454402 247052 454408 247064
rect 454460 247052 454466 247104
rect 443638 245556 443644 245608
rect 443696 245596 443702 245608
rect 580166 245596 580172 245608
rect 443696 245568 580172 245596
rect 443696 245556 443702 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 442902 244264 442908 244316
rect 442960 244304 442966 244316
rect 451550 244304 451556 244316
rect 442960 244276 451556 244304
rect 442960 244264 442966 244276
rect 451550 244264 451556 244276
rect 451608 244264 451614 244316
rect 51166 242904 51172 242956
rect 51224 242944 51230 242956
rect 57330 242944 57336 242956
rect 51224 242916 57336 242944
rect 51224 242904 51230 242916
rect 57330 242904 57336 242916
rect 57388 242904 57394 242956
rect 3050 241408 3056 241460
rect 3108 241448 3114 241460
rect 54294 241448 54300 241460
rect 3108 241420 54300 241448
rect 3108 241408 3114 241420
rect 54294 241408 54300 241420
rect 54352 241408 54358 241460
rect 442718 239096 442724 239148
rect 442776 239136 442782 239148
rect 443822 239136 443828 239148
rect 442776 239108 443828 239136
rect 442776 239096 442782 239108
rect 443822 239096 443828 239108
rect 443880 239096 443886 239148
rect 46566 238756 46572 238808
rect 46624 238796 46630 238808
rect 57330 238796 57336 238808
rect 46624 238768 57336 238796
rect 46624 238756 46630 238768
rect 57330 238756 57336 238768
rect 57388 238756 57394 238808
rect 442902 235968 442908 236020
rect 442960 236008 442966 236020
rect 453022 236008 453028 236020
rect 442960 235980 453028 236008
rect 442960 235968 442966 235980
rect 453022 235968 453028 235980
rect 453080 235968 453086 236020
rect 442902 233384 442908 233436
rect 442960 233424 442966 233436
rect 445754 233424 445760 233436
rect 442960 233396 445760 233424
rect 442960 233384 442966 233396
rect 445754 233384 445760 233396
rect 445812 233384 445818 233436
rect 442902 230664 442908 230716
rect 442960 230704 442966 230716
rect 449158 230704 449164 230716
rect 442960 230676 449164 230704
rect 442960 230664 442966 230676
rect 449158 230664 449164 230676
rect 449216 230664 449222 230716
rect 54294 230460 54300 230512
rect 54352 230500 54358 230512
rect 57330 230500 57336 230512
rect 54352 230472 57336 230500
rect 54352 230460 54358 230472
rect 57330 230460 57336 230472
rect 57388 230460 57394 230512
rect 57330 230324 57336 230376
rect 57388 230364 57394 230376
rect 57882 230364 57888 230376
rect 57388 230336 57888 230364
rect 57388 230324 57394 230336
rect 57882 230324 57888 230336
rect 57940 230324 57946 230376
rect 50338 227740 50344 227792
rect 50396 227780 50402 227792
rect 57882 227780 57888 227792
rect 50396 227752 57888 227780
rect 50396 227740 50402 227752
rect 57882 227740 57888 227752
rect 57940 227740 57946 227792
rect 442902 226312 442908 226364
rect 442960 226352 442966 226364
rect 480254 226352 480260 226364
rect 442960 226324 480260 226352
rect 442960 226312 442966 226324
rect 480254 226312 480260 226324
rect 480312 226312 480318 226364
rect 52546 224952 52552 225004
rect 52604 224992 52610 225004
rect 57882 224992 57888 225004
rect 52604 224964 57888 224992
rect 52604 224952 52610 224964
rect 57882 224952 57888 224964
rect 57940 224952 57946 225004
rect 45094 222164 45100 222216
rect 45152 222204 45158 222216
rect 57882 222204 57888 222216
rect 45152 222176 57888 222204
rect 45152 222164 45158 222176
rect 57882 222164 57888 222176
rect 57940 222164 57946 222216
rect 442626 221008 442632 221060
rect 442684 221048 442690 221060
rect 443638 221048 443644 221060
rect 442684 221020 443644 221048
rect 442684 221008 442690 221020
rect 443638 221008 443644 221020
rect 443696 221008 443702 221060
rect 508498 219376 508504 219428
rect 508556 219416 508562 219428
rect 579982 219416 579988 219428
rect 508556 219388 579988 219416
rect 508556 219376 508562 219388
rect 579982 219376 579988 219388
rect 580040 219376 580046 219428
rect 54110 218016 54116 218068
rect 54168 218056 54174 218068
rect 57882 218056 57888 218068
rect 54168 218028 57888 218056
rect 54168 218016 54174 218028
rect 57882 218016 57888 218028
rect 57940 218016 57946 218068
rect 442902 218016 442908 218068
rect 442960 218056 442966 218068
rect 507854 218056 507860 218068
rect 442960 218028 507860 218056
rect 442960 218016 442966 218028
rect 507854 218016 507860 218028
rect 507912 218016 507918 218068
rect 55766 215296 55772 215348
rect 55824 215336 55830 215348
rect 56594 215336 56600 215348
rect 55824 215308 56600 215336
rect 55824 215296 55830 215308
rect 56594 215296 56600 215308
rect 56652 215296 56658 215348
rect 442902 215296 442908 215348
rect 442960 215336 442966 215348
rect 545758 215336 545764 215348
rect 442960 215308 545764 215336
rect 442960 215296 442966 215308
rect 545758 215296 545764 215308
rect 545816 215296 545822 215348
rect 442718 212848 442724 212900
rect 442776 212888 442782 212900
rect 444006 212888 444012 212900
rect 442776 212860 444012 212888
rect 442776 212848 442782 212860
rect 444006 212848 444012 212860
rect 444064 212848 444070 212900
rect 442718 210264 442724 210316
rect 442776 210304 442782 210316
rect 450446 210304 450452 210316
rect 442776 210276 450452 210304
rect 442776 210264 442782 210276
rect 450446 210264 450452 210276
rect 450504 210264 450510 210316
rect 3510 209788 3516 209840
rect 3568 209828 3574 209840
rect 57882 209828 57888 209840
rect 3568 209800 57888 209828
rect 3568 209788 3574 209800
rect 57882 209788 57888 209800
rect 57940 209788 57946 209840
rect 57790 208496 57796 208548
rect 57848 208496 57854 208548
rect 57808 208344 57836 208496
rect 49510 208292 49516 208344
rect 49568 208332 49574 208344
rect 57698 208332 57704 208344
rect 49568 208304 57704 208332
rect 49568 208292 49574 208304
rect 57698 208292 57704 208304
rect 57756 208292 57762 208344
rect 57790 208292 57796 208344
rect 57848 208292 57854 208344
rect 53926 204280 53932 204332
rect 53984 204320 53990 204332
rect 57698 204320 57704 204332
rect 53984 204292 57704 204320
rect 53984 204280 53990 204292
rect 57698 204280 57704 204292
rect 57756 204280 57762 204332
rect 442902 204212 442908 204264
rect 442960 204252 442966 204264
rect 464338 204252 464344 204264
rect 442960 204224 464344 204252
rect 442960 204212 442966 204224
rect 464338 204212 464344 204224
rect 464396 204212 464402 204264
rect 442902 201492 442908 201544
rect 442960 201532 442966 201544
rect 537478 201532 537484 201544
rect 442960 201504 537484 201532
rect 442960 201492 442966 201504
rect 537478 201492 537484 201504
rect 537536 201492 537542 201544
rect 55582 198704 55588 198756
rect 55640 198744 55646 198756
rect 56594 198744 56600 198756
rect 55640 198716 56600 198744
rect 55640 198704 55646 198716
rect 56594 198704 56600 198716
rect 56652 198704 56658 198756
rect 442902 198704 442908 198756
rect 442960 198744 442966 198756
rect 453114 198744 453120 198756
rect 442960 198716 453120 198744
rect 442960 198704 442966 198716
rect 453114 198704 453120 198716
rect 453172 198704 453178 198756
rect 44910 195984 44916 196036
rect 44968 196024 44974 196036
rect 57698 196024 57704 196036
rect 44968 195996 57704 196024
rect 44968 195984 44974 195996
rect 57698 195984 57704 195996
rect 57756 195984 57762 196036
rect 442902 195304 442908 195356
rect 442960 195344 442966 195356
rect 444742 195344 444748 195356
rect 442960 195316 444748 195344
rect 442960 195304 442966 195316
rect 444742 195304 444748 195316
rect 444800 195304 444806 195356
rect 45370 194488 45376 194540
rect 45428 194528 45434 194540
rect 57698 194528 57704 194540
rect 45428 194500 57704 194528
rect 45428 194488 45434 194500
rect 57698 194488 57704 194500
rect 57756 194488 57762 194540
rect 442902 192584 442908 192636
rect 442960 192624 442966 192636
rect 450538 192624 450544 192636
rect 442960 192596 450544 192624
rect 442960 192584 442966 192596
rect 450538 192584 450544 192596
rect 450596 192584 450602 192636
rect 53834 190476 53840 190528
rect 53892 190516 53898 190528
rect 56870 190516 56876 190528
rect 53892 190488 56876 190516
rect 53892 190476 53898 190488
rect 56870 190476 56876 190488
rect 56928 190476 56934 190528
rect 3326 188980 3332 189032
rect 3384 189020 3390 189032
rect 18598 189020 18604 189032
rect 3384 188992 18604 189020
rect 3384 188980 3390 188992
rect 18598 188980 18604 188992
rect 18656 188980 18662 189032
rect 3234 187620 3240 187672
rect 3292 187660 3298 187672
rect 57698 187660 57704 187672
rect 3292 187632 57704 187660
rect 3292 187620 3298 187632
rect 57698 187620 57704 187632
rect 57756 187620 57762 187672
rect 442626 186464 442632 186516
rect 442684 186504 442690 186516
rect 443730 186504 443736 186516
rect 442684 186476 443736 186504
rect 442684 186464 442690 186476
rect 443730 186464 443736 186476
rect 443788 186464 443794 186516
rect 46474 183540 46480 183592
rect 46532 183580 46538 183592
rect 57698 183580 57704 183592
rect 46532 183552 57704 183580
rect 46532 183540 46538 183552
rect 57698 183540 57704 183552
rect 57756 183540 57762 183592
rect 442902 181024 442908 181076
rect 442960 181064 442966 181076
rect 446490 181064 446496 181076
rect 442960 181036 446496 181064
rect 442960 181024 442966 181036
rect 446490 181024 446496 181036
rect 446548 181024 446554 181076
rect 3970 180820 3976 180872
rect 4028 180860 4034 180872
rect 57698 180860 57704 180872
rect 4028 180832 57704 180860
rect 4028 180820 4034 180832
rect 57698 180820 57704 180832
rect 57756 180820 57762 180872
rect 442902 178304 442908 178356
rect 442960 178344 442966 178356
rect 450630 178344 450636 178356
rect 442960 178316 450636 178344
rect 442960 178304 442966 178316
rect 450630 178304 450636 178316
rect 450688 178304 450694 178356
rect 442718 175584 442724 175636
rect 442776 175624 442782 175636
rect 444834 175624 444840 175636
rect 442776 175596 444840 175624
rect 442776 175584 442782 175596
rect 444834 175584 444840 175596
rect 444892 175584 444898 175636
rect 49510 172524 49516 172576
rect 49568 172564 49574 172576
rect 57698 172564 57704 172576
rect 49568 172536 57704 172564
rect 49568 172524 49574 172536
rect 57698 172524 57704 172536
rect 57756 172524 57762 172576
rect 57790 172456 57796 172508
rect 57848 172456 57854 172508
rect 57808 172304 57836 172456
rect 57790 172252 57796 172304
rect 57848 172252 57854 172304
rect 442902 171096 442908 171148
rect 442960 171136 442966 171148
rect 525794 171136 525800 171148
rect 442960 171108 525800 171136
rect 442960 171096 442966 171108
rect 525794 171096 525800 171108
rect 525852 171096 525858 171148
rect 41322 171028 41328 171080
rect 41380 171068 41386 171080
rect 57882 171068 57888 171080
rect 41380 171040 57888 171068
rect 41380 171028 41386 171040
rect 57882 171028 57888 171040
rect 57940 171028 57946 171080
rect 442902 168376 442908 168428
rect 442960 168416 442966 168428
rect 451642 168416 451648 168428
rect 442960 168388 451648 168416
rect 442960 168376 442966 168388
rect 451642 168376 451648 168388
rect 451700 168376 451706 168428
rect 47670 165588 47676 165640
rect 47728 165628 47734 165640
rect 57882 165628 57888 165640
rect 47728 165600 57888 165628
rect 47728 165588 47734 165600
rect 57882 165588 57888 165600
rect 57940 165588 57946 165640
rect 49326 162868 49332 162920
rect 49384 162908 49390 162920
rect 57882 162908 57888 162920
rect 49384 162880 57888 162908
rect 49384 162868 49390 162880
rect 57882 162868 57888 162880
rect 57940 162868 57946 162920
rect 442902 160624 442908 160676
rect 442960 160664 442966 160676
rect 444926 160664 444932 160676
rect 442960 160636 444932 160664
rect 442960 160624 442966 160636
rect 444926 160624 444932 160636
rect 444984 160624 444990 160676
rect 442718 158652 442724 158704
rect 442776 158692 442782 158704
rect 580810 158692 580816 158704
rect 442776 158664 580816 158692
rect 442776 158652 442782 158664
rect 580810 158652 580816 158664
rect 580868 158652 580874 158704
rect 47946 155864 47952 155916
rect 48004 155904 48010 155916
rect 57882 155904 57888 155916
rect 48004 155876 57888 155904
rect 48004 155864 48010 155876
rect 57882 155864 57888 155876
rect 57940 155864 57946 155916
rect 439498 152464 439504 152516
rect 439556 152464 439562 152516
rect 439590 152464 439596 152516
rect 439648 152464 439654 152516
rect 439516 152312 439544 152464
rect 439608 152312 439636 152464
rect 439498 152260 439504 152312
rect 439556 152260 439562 152312
rect 439590 152260 439596 152312
rect 439648 152260 439654 152312
rect 26142 151784 26148 151836
rect 26200 151824 26206 151836
rect 57882 151824 57888 151836
rect 26200 151796 57888 151824
rect 26200 151784 26206 151796
rect 57882 151784 57888 151796
rect 57940 151784 57946 151836
rect 2774 150084 2780 150136
rect 2832 150124 2838 150136
rect 4798 150124 4804 150136
rect 2832 150096 4804 150124
rect 2832 150084 2838 150096
rect 4798 150084 4804 150096
rect 4856 150084 4862 150136
rect 51074 149200 51080 149252
rect 51132 149240 51138 149252
rect 54202 149240 54208 149252
rect 51132 149212 54208 149240
rect 51132 149200 51138 149212
rect 54202 149200 54208 149212
rect 54260 149200 54266 149252
rect 54202 149064 54208 149116
rect 54260 149104 54266 149116
rect 57882 149104 57888 149116
rect 54260 149076 57888 149104
rect 54260 149064 54266 149076
rect 57882 149064 57888 149076
rect 57940 149064 57946 149116
rect 442902 149064 442908 149116
rect 442960 149104 442966 149116
rect 500954 149104 500960 149116
rect 442960 149076 500960 149104
rect 442960 149064 442966 149076
rect 500954 149064 500960 149076
rect 501012 149064 501018 149116
rect 442810 147568 442816 147620
rect 442868 147608 442874 147620
rect 580902 147608 580908 147620
rect 442868 147580 580908 147608
rect 442868 147568 442874 147580
rect 580902 147568 580908 147580
rect 580960 147568 580966 147620
rect 52454 146616 52460 146668
rect 52512 146656 52518 146668
rect 54018 146656 54024 146668
rect 52512 146628 54024 146656
rect 52512 146616 52518 146628
rect 54018 146616 54024 146628
rect 54076 146616 54082 146668
rect 54018 146276 54024 146328
rect 54076 146316 54082 146328
rect 57882 146316 57888 146328
rect 54076 146288 57888 146316
rect 54076 146276 54082 146288
rect 57882 146276 57888 146288
rect 57940 146276 57946 146328
rect 442902 143624 442908 143676
rect 442960 143664 442966 143676
rect 449250 143664 449256 143676
rect 442960 143636 449256 143664
rect 442960 143624 442966 143636
rect 449250 143624 449256 143636
rect 449308 143624 449314 143676
rect 46290 140768 46296 140820
rect 46348 140808 46354 140820
rect 57882 140808 57888 140820
rect 46348 140780 57888 140808
rect 46348 140768 46354 140780
rect 57882 140768 57888 140780
rect 57940 140768 57946 140820
rect 442902 139408 442908 139460
rect 442960 139448 442966 139460
rect 460198 139448 460204 139460
rect 442960 139420 460204 139448
rect 442960 139408 442966 139420
rect 460198 139408 460204 139420
rect 460256 139408 460262 139460
rect 3326 137912 3332 137964
rect 3384 137952 3390 137964
rect 29638 137952 29644 137964
rect 3384 137924 29644 137952
rect 3384 137912 3390 137924
rect 29638 137912 29644 137924
rect 29696 137912 29702 137964
rect 47946 135260 47952 135312
rect 48004 135300 48010 135312
rect 57882 135300 57888 135312
rect 48004 135272 57888 135300
rect 48004 135260 48010 135272
rect 57882 135260 57888 135272
rect 57940 135260 57946 135312
rect 442902 132064 442908 132116
rect 442960 132104 442966 132116
rect 446582 132104 446588 132116
rect 442960 132076 446588 132104
rect 442960 132064 442966 132076
rect 446582 132064 446588 132076
rect 446640 132064 446646 132116
rect 47578 131112 47584 131164
rect 47636 131152 47642 131164
rect 57882 131152 57888 131164
rect 47636 131124 57888 131152
rect 47636 131112 47642 131124
rect 57882 131112 57888 131124
rect 57940 131112 57946 131164
rect 49234 128324 49240 128376
rect 49292 128364 49298 128376
rect 57882 128364 57888 128376
rect 49292 128336 57888 128364
rect 49292 128324 49298 128336
rect 57882 128324 57888 128336
rect 57940 128324 57946 128376
rect 441522 125604 441528 125656
rect 441580 125644 441586 125656
rect 465074 125644 465080 125656
rect 441580 125616 465080 125644
rect 441580 125604 441586 125616
rect 465074 125604 465080 125616
rect 465132 125604 465138 125656
rect 46382 122816 46388 122868
rect 46440 122856 46446 122868
rect 57882 122856 57888 122868
rect 46440 122828 57888 122856
rect 46440 122816 46446 122828
rect 57882 122816 57888 122828
rect 57940 122816 57946 122868
rect 441522 122816 441528 122868
rect 441580 122856 441586 122868
rect 446766 122856 446772 122868
rect 441580 122828 446772 122856
rect 441580 122816 441586 122828
rect 446766 122816 446772 122828
rect 446824 122816 446830 122868
rect 50246 120096 50252 120148
rect 50304 120136 50310 120148
rect 57882 120136 57888 120148
rect 50304 120108 57888 120136
rect 50304 120096 50310 120108
rect 57882 120096 57888 120108
rect 57940 120096 57946 120148
rect 441522 118668 441528 118720
rect 441580 118708 441586 118720
rect 445018 118708 445024 118720
rect 441580 118680 445024 118708
rect 441580 118668 441586 118680
rect 445018 118668 445024 118680
rect 445076 118668 445082 118720
rect 49142 117308 49148 117360
rect 49200 117348 49206 117360
rect 57882 117348 57888 117360
rect 49200 117320 57888 117348
rect 49200 117308 49206 117320
rect 57882 117308 57888 117320
rect 57940 117308 57946 117360
rect 441522 115948 441528 116000
rect 441580 115988 441586 116000
rect 494698 115988 494704 116000
rect 441580 115960 494704 115988
rect 441580 115948 441586 115960
rect 494698 115948 494704 115960
rect 494756 115948 494762 116000
rect 47486 114520 47492 114572
rect 47544 114560 47550 114572
rect 57882 114560 57888 114572
rect 47544 114532 57888 114560
rect 47544 114520 47550 114532
rect 57882 114520 57888 114532
rect 57940 114520 57946 114572
rect 441522 114384 441528 114436
rect 441580 114424 441586 114436
rect 444098 114424 444104 114436
rect 441580 114396 444104 114424
rect 441580 114384 441586 114396
rect 444098 114384 444104 114396
rect 444156 114384 444162 114436
rect 454678 113092 454684 113144
rect 454736 113132 454742 113144
rect 579982 113132 579988 113144
rect 454736 113104 579988 113132
rect 454736 113092 454742 113104
rect 579982 113092 579988 113104
rect 580040 113092 580046 113144
rect 441522 110440 441528 110492
rect 441580 110480 441586 110492
rect 451458 110480 451464 110492
rect 441580 110452 451464 110480
rect 441580 110440 441586 110452
rect 451458 110440 451464 110452
rect 451516 110440 451522 110492
rect 441522 107652 441528 107704
rect 441580 107692 441586 107704
rect 515398 107692 515404 107704
rect 441580 107664 515404 107692
rect 441580 107652 441586 107664
rect 515398 107652 515404 107664
rect 515456 107652 515462 107704
rect 48222 107584 48228 107636
rect 48280 107624 48286 107636
rect 57882 107624 57888 107636
rect 48280 107596 57888 107624
rect 48280 107584 48286 107596
rect 57882 107584 57888 107596
rect 57940 107584 57946 107636
rect 441522 104864 441528 104916
rect 441580 104904 441586 104916
rect 477494 104904 477500 104916
rect 441580 104876 477500 104904
rect 441580 104864 441586 104876
rect 477494 104864 477500 104876
rect 477552 104864 477558 104916
rect 55490 103504 55496 103556
rect 55548 103544 55554 103556
rect 56594 103544 56600 103556
rect 55548 103516 56600 103544
rect 55548 103504 55554 103516
rect 56594 103504 56600 103516
rect 56652 103504 56658 103556
rect 441522 103436 441528 103488
rect 441580 103476 441586 103488
rect 446030 103476 446036 103488
rect 441580 103448 446036 103476
rect 441580 103436 441586 103448
rect 446030 103436 446036 103448
rect 446088 103436 446094 103488
rect 48038 100648 48044 100700
rect 48096 100688 48102 100700
rect 57882 100688 57888 100700
rect 48096 100660 57888 100688
rect 48096 100648 48102 100660
rect 57882 100648 57888 100660
rect 57940 100648 57946 100700
rect 566458 100648 566464 100700
rect 566516 100688 566522 100700
rect 580166 100688 580172 100700
rect 566516 100660 580172 100688
rect 566516 100648 566522 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 441522 99356 441528 99408
rect 441580 99396 441586 99408
rect 446674 99396 446680 99408
rect 441580 99368 446680 99396
rect 441580 99356 441586 99368
rect 446674 99356 446680 99368
rect 446732 99356 446738 99408
rect 50154 93848 50160 93900
rect 50212 93888 50218 93900
rect 57882 93888 57888 93900
rect 50212 93860 57888 93888
rect 50212 93848 50218 93860
rect 57882 93848 57888 93860
rect 57940 93848 57946 93900
rect 441522 91060 441528 91112
rect 441580 91100 441586 91112
rect 461670 91100 461676 91112
rect 441580 91072 461676 91100
rect 441580 91060 441586 91072
rect 461670 91060 461676 91072
rect 461728 91060 461734 91112
rect 443914 88000 443920 88052
rect 443972 88040 443978 88052
rect 445018 88040 445024 88052
rect 443972 88012 445024 88040
rect 443972 88000 443978 88012
rect 445018 88000 445024 88012
rect 445076 88000 445082 88052
rect 441522 86980 441528 87032
rect 441580 87020 441586 87032
rect 548518 87020 548524 87032
rect 441580 86992 548524 87020
rect 441580 86980 441586 86992
rect 548518 86980 548524 86992
rect 548576 86980 548582 87032
rect 57882 86000 57888 86012
rect 57843 85972 57888 86000
rect 57882 85960 57888 85972
rect 57940 85960 57946 86012
rect 33042 85552 33048 85604
rect 33100 85592 33106 85604
rect 57882 85592 57888 85604
rect 33100 85564 57888 85592
rect 33100 85552 33106 85564
rect 57882 85552 57888 85564
rect 57940 85552 57946 85604
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 21358 85524 21364 85536
rect 3384 85496 21364 85524
rect 3384 85484 3390 85496
rect 21358 85484 21364 85496
rect 21416 85484 21422 85536
rect 57882 85456 57888 85468
rect 57843 85428 57888 85456
rect 57882 85416 57888 85428
rect 57940 85416 57946 85468
rect 441522 81404 441528 81456
rect 441580 81444 441586 81456
rect 445018 81444 445024 81456
rect 441580 81416 445024 81444
rect 441580 81404 441586 81416
rect 445018 81404 445024 81416
rect 445076 81404 445082 81456
rect 441522 79976 441528 80028
rect 441580 80016 441586 80028
rect 449894 80016 449900 80028
rect 441580 79988 449900 80016
rect 441580 79976 441586 79988
rect 449894 79976 449900 79988
rect 449952 79976 449958 80028
rect 14458 77188 14464 77240
rect 14516 77228 14522 77240
rect 56870 77228 56876 77240
rect 14516 77200 56876 77228
rect 14516 77188 14522 77200
rect 56870 77188 56876 77200
rect 56928 77188 56934 77240
rect 441522 76304 441528 76356
rect 441580 76344 441586 76356
rect 445110 76344 445116 76356
rect 441580 76316 445116 76344
rect 441580 76304 441586 76316
rect 445110 76304 445116 76316
rect 445168 76304 445174 76356
rect 439498 73176 439504 73228
rect 439556 73176 439562 73228
rect 439516 73024 439544 73176
rect 439498 72972 439504 73024
rect 439556 72972 439562 73024
rect 3510 68416 3516 68468
rect 3568 68456 3574 68468
rect 3694 68456 3700 68468
rect 3568 68428 3700 68456
rect 3568 68416 3574 68428
rect 3694 68416 3700 68428
rect 3752 68416 3758 68468
rect 17218 66172 17224 66224
rect 17276 66212 17282 66224
rect 56870 66212 56876 66224
rect 17276 66184 56876 66212
rect 17276 66172 17282 66184
rect 56870 66172 56876 66184
rect 56928 66172 56934 66224
rect 58066 61752 58072 61804
rect 58124 61792 58130 61804
rect 302237 61795 302295 61801
rect 302237 61792 302249 61795
rect 58124 61764 302249 61792
rect 58124 61752 58130 61764
rect 302237 61761 302249 61764
rect 302283 61761 302295 61795
rect 302237 61755 302295 61761
rect 315945 61795 316003 61801
rect 315945 61761 315957 61795
rect 315991 61792 316003 61795
rect 443546 61792 443552 61804
rect 315991 61764 443552 61792
rect 315991 61761 316003 61764
rect 315945 61755 316003 61761
rect 443546 61752 443552 61764
rect 443604 61752 443610 61804
rect 58986 61684 58992 61736
rect 59044 61724 59050 61736
rect 358817 61727 358875 61733
rect 358817 61724 358829 61727
rect 59044 61696 358829 61724
rect 59044 61684 59050 61696
rect 358817 61693 358829 61696
rect 358863 61693 358875 61727
rect 358817 61687 358875 61693
rect 375285 61727 375343 61733
rect 375285 61693 375297 61727
rect 375331 61724 375343 61727
rect 444006 61724 444012 61736
rect 375331 61696 444012 61724
rect 375331 61693 375343 61696
rect 375285 61687 375343 61693
rect 444006 61684 444012 61696
rect 444064 61684 444070 61736
rect 52086 61616 52092 61668
rect 52144 61656 52150 61668
rect 375377 61659 375435 61665
rect 375377 61656 375389 61659
rect 52144 61628 375389 61656
rect 52144 61616 52150 61628
rect 375377 61625 375389 61628
rect 375423 61625 375435 61659
rect 375377 61619 375435 61625
rect 378045 61659 378103 61665
rect 378045 61625 378057 61659
rect 378091 61656 378103 61659
rect 441246 61656 441252 61668
rect 378091 61628 441252 61656
rect 378091 61625 378103 61628
rect 378045 61619 378103 61625
rect 441246 61616 441252 61628
rect 441304 61616 441310 61668
rect 56318 61548 56324 61600
rect 56376 61588 56382 61600
rect 484394 61588 484400 61600
rect 56376 61560 484400 61588
rect 56376 61548 56382 61560
rect 484394 61548 484400 61560
rect 484452 61548 484458 61600
rect 58434 61480 58440 61532
rect 58492 61520 58498 61532
rect 488534 61520 488540 61532
rect 58492 61492 488540 61520
rect 58492 61480 58498 61492
rect 488534 61480 488540 61492
rect 488592 61480 488598 61532
rect 55582 61412 55588 61464
rect 55640 61452 55646 61464
rect 498286 61452 498292 61464
rect 55640 61424 498292 61452
rect 55640 61412 55646 61424
rect 498286 61412 498292 61424
rect 498344 61412 498350 61464
rect 56226 61344 56232 61396
rect 56284 61384 56290 61396
rect 509234 61384 509240 61396
rect 56284 61356 509240 61384
rect 56284 61344 56290 61356
rect 509234 61344 509240 61356
rect 509292 61344 509298 61396
rect 58618 61276 58624 61328
rect 58676 61316 58682 61328
rect 168377 61319 168435 61325
rect 168377 61316 168389 61319
rect 58676 61288 168389 61316
rect 58676 61276 58682 61288
rect 168377 61285 168389 61288
rect 168423 61285 168435 61319
rect 168377 61279 168435 61285
rect 211065 61319 211123 61325
rect 211065 61285 211077 61319
rect 211111 61316 211123 61319
rect 441154 61316 441160 61328
rect 211111 61288 441160 61316
rect 211111 61285 211123 61288
rect 211065 61279 211123 61285
rect 441154 61276 441160 61288
rect 441212 61276 441218 61328
rect 54018 61208 54024 61260
rect 54076 61248 54082 61260
rect 218057 61251 218115 61257
rect 218057 61248 218069 61251
rect 54076 61220 218069 61248
rect 54076 61208 54082 61220
rect 218057 61217 218069 61220
rect 218103 61217 218115 61251
rect 218057 61211 218115 61217
rect 224681 61251 224739 61257
rect 224681 61217 224693 61251
rect 224727 61248 224739 61251
rect 446306 61248 446312 61260
rect 224727 61220 446312 61248
rect 224727 61217 224739 61220
rect 224681 61211 224739 61217
rect 446306 61208 446312 61220
rect 446364 61208 446370 61260
rect 55674 61140 55680 61192
rect 55732 61180 55738 61192
rect 258077 61183 258135 61189
rect 258077 61180 258089 61183
rect 55732 61152 258089 61180
rect 55732 61140 55738 61152
rect 258077 61149 258089 61152
rect 258123 61149 258135 61183
rect 258077 61143 258135 61149
rect 286965 61183 287023 61189
rect 286965 61149 286977 61183
rect 287011 61180 287023 61183
rect 444098 61180 444104 61192
rect 287011 61152 444104 61180
rect 287011 61149 287023 61152
rect 286965 61143 287023 61149
rect 444098 61140 444104 61152
rect 444156 61140 444162 61192
rect 54478 61072 54484 61124
rect 54536 61112 54542 61124
rect 254029 61115 254087 61121
rect 254029 61112 254041 61115
rect 54536 61084 254041 61112
rect 54536 61072 54542 61084
rect 254029 61081 254041 61084
rect 254075 61081 254087 61115
rect 254029 61075 254087 61081
rect 257985 61115 258043 61121
rect 257985 61081 257997 61115
rect 258031 61112 258043 61115
rect 440510 61112 440516 61124
rect 258031 61084 440516 61112
rect 258031 61081 258043 61084
rect 257985 61075 258043 61081
rect 440510 61072 440516 61084
rect 440568 61072 440574 61124
rect 53834 61004 53840 61056
rect 53892 61044 53898 61056
rect 235997 61047 236055 61053
rect 235997 61044 236009 61047
rect 53892 61016 236009 61044
rect 53892 61004 53898 61016
rect 235997 61013 236009 61016
rect 236043 61013 236055 61047
rect 235997 61007 236055 61013
rect 291105 61047 291163 61053
rect 291105 61013 291117 61047
rect 291151 61044 291163 61047
rect 439682 61044 439688 61056
rect 291151 61016 439688 61044
rect 291151 61013 291163 61016
rect 291105 61007 291163 61013
rect 439682 61004 439688 61016
rect 439740 61004 439746 61056
rect 51534 60936 51540 60988
rect 51592 60976 51598 60988
rect 149149 60979 149207 60985
rect 149149 60976 149161 60979
rect 51592 60948 149161 60976
rect 51592 60936 51598 60948
rect 149149 60945 149161 60948
rect 149195 60945 149207 60979
rect 149149 60939 149207 60945
rect 350445 60979 350503 60985
rect 350445 60945 350457 60979
rect 350491 60976 350503 60979
rect 444650 60976 444656 60988
rect 350491 60948 444656 60976
rect 350491 60945 350503 60948
rect 350445 60939 350503 60945
rect 444650 60936 444656 60948
rect 444708 60936 444714 60988
rect 58526 60868 58532 60920
rect 58584 60908 58590 60920
rect 143537 60911 143595 60917
rect 143537 60908 143549 60911
rect 58584 60880 143549 60908
rect 58584 60868 58590 60880
rect 143537 60877 143549 60880
rect 143583 60877 143595 60911
rect 143537 60871 143595 60877
rect 400125 60911 400183 60917
rect 400125 60877 400137 60911
rect 400171 60908 400183 60911
rect 440786 60908 440792 60920
rect 400171 60880 440792 60908
rect 400171 60877 400183 60880
rect 400125 60871 400183 60877
rect 440786 60868 440792 60880
rect 440844 60868 440850 60920
rect 441522 60868 441528 60920
rect 441580 60908 441586 60920
rect 507118 60908 507124 60920
rect 441580 60880 507124 60908
rect 441580 60868 441586 60880
rect 507118 60868 507124 60880
rect 507176 60868 507182 60920
rect 54662 60800 54668 60852
rect 54720 60840 54726 60852
rect 80057 60843 80115 60849
rect 80057 60840 80069 60843
rect 54720 60812 80069 60840
rect 54720 60800 54726 60812
rect 80057 60809 80069 60812
rect 80103 60809 80115 60843
rect 80057 60803 80115 60809
rect 404265 60843 404323 60849
rect 404265 60809 404277 60843
rect 404311 60840 404323 60843
rect 444834 60840 444840 60852
rect 404311 60812 444840 60840
rect 404311 60809 404323 60812
rect 404265 60803 404323 60809
rect 444834 60800 444840 60812
rect 444892 60800 444898 60852
rect 431865 60775 431923 60781
rect 431865 60741 431877 60775
rect 431911 60772 431923 60775
rect 443178 60772 443184 60784
rect 431911 60744 443184 60772
rect 431911 60741 431923 60744
rect 431865 60735 431923 60741
rect 443178 60732 443184 60744
rect 443236 60732 443242 60784
rect 46658 60664 46664 60716
rect 46716 60704 46722 60716
rect 580534 60704 580540 60716
rect 46716 60676 580540 60704
rect 46716 60664 46722 60676
rect 580534 60664 580540 60676
rect 580592 60664 580598 60716
rect 50246 60596 50252 60648
rect 50304 60636 50310 60648
rect 176654 60636 176660 60648
rect 50304 60608 176660 60636
rect 50304 60596 50310 60608
rect 176654 60596 176660 60608
rect 176712 60596 176718 60648
rect 200022 60596 200028 60648
rect 200080 60636 200086 60648
rect 445938 60636 445944 60648
rect 200080 60608 445944 60636
rect 200080 60596 200086 60608
rect 445938 60596 445944 60608
rect 445996 60596 446002 60648
rect 49602 60528 49608 60580
rect 49660 60568 49666 60580
rect 160094 60568 160100 60580
rect 49660 60540 160100 60568
rect 49660 60528 49666 60540
rect 160094 60528 160100 60540
rect 160152 60528 160158 60580
rect 168282 60528 168288 60580
rect 168340 60568 168346 60580
rect 444558 60568 444564 60580
rect 168340 60540 444564 60568
rect 168340 60528 168346 60540
rect 444558 60528 444564 60540
rect 444616 60528 444622 60580
rect 51994 60460 52000 60512
rect 52052 60500 52058 60512
rect 336734 60500 336740 60512
rect 52052 60472 336740 60500
rect 52052 60460 52058 60472
rect 336734 60460 336740 60472
rect 336792 60460 336798 60512
rect 350442 60500 350448 60512
rect 350403 60472 350448 60500
rect 350442 60460 350448 60472
rect 350500 60460 350506 60512
rect 358722 60460 358728 60512
rect 358780 60500 358786 60512
rect 444926 60500 444932 60512
rect 358780 60472 444932 60500
rect 358780 60460 358786 60472
rect 444926 60460 444932 60472
rect 444984 60460 444990 60512
rect 59906 60392 59912 60444
rect 59964 60432 59970 60444
rect 135254 60432 135260 60444
rect 59964 60404 135260 60432
rect 59964 60392 59970 60404
rect 135254 60392 135260 60404
rect 135312 60392 135318 60444
rect 143534 60432 143540 60444
rect 143495 60404 143540 60432
rect 143534 60392 143540 60404
rect 143592 60392 143598 60444
rect 149146 60432 149152 60444
rect 149107 60404 149152 60432
rect 149146 60392 149152 60404
rect 149204 60392 149210 60444
rect 151722 60392 151728 60444
rect 151780 60432 151786 60444
rect 443822 60432 443828 60444
rect 151780 60404 443828 60432
rect 151780 60392 151786 60404
rect 443822 60392 443828 60404
rect 443880 60392 443886 60444
rect 59262 60324 59268 60376
rect 59320 60364 59326 60376
rect 67634 60364 67640 60376
rect 59320 60336 67640 60364
rect 59320 60324 59326 60336
rect 67634 60324 67640 60336
rect 67692 60324 67698 60376
rect 80054 60364 80060 60376
rect 80015 60336 80060 60364
rect 80054 60324 80060 60336
rect 80112 60324 80118 60376
rect 122742 60324 122748 60376
rect 122800 60364 122806 60376
rect 447962 60364 447968 60376
rect 122800 60336 447968 60364
rect 122800 60324 122806 60336
rect 447962 60324 447968 60336
rect 448020 60324 448026 60376
rect 56686 60256 56692 60308
rect 56744 60296 56750 60308
rect 82814 60296 82820 60308
rect 56744 60268 82820 60296
rect 56744 60256 56750 60268
rect 82814 60256 82820 60268
rect 82872 60256 82878 60308
rect 99282 60256 99288 60308
rect 99340 60296 99346 60308
rect 448238 60296 448244 60308
rect 99340 60268 448244 60296
rect 99340 60256 99346 60268
rect 448238 60256 448244 60268
rect 448296 60256 448302 60308
rect 45002 60188 45008 60240
rect 45060 60228 45066 60240
rect 448146 60228 448152 60240
rect 45060 60200 448152 60228
rect 45060 60188 45066 60200
rect 448146 60188 448152 60200
rect 448204 60188 448210 60240
rect 6822 60120 6828 60172
rect 6880 60160 6886 60172
rect 449066 60160 449072 60172
rect 6880 60132 449072 60160
rect 6880 60120 6886 60132
rect 449066 60120 449072 60132
rect 449124 60120 449130 60172
rect 52638 60052 52644 60104
rect 52696 60092 52702 60104
rect 549254 60092 549260 60104
rect 52696 60064 549260 60092
rect 52696 60052 52702 60064
rect 549254 60052 549260 60064
rect 549312 60052 549318 60104
rect 52822 59984 52828 60036
rect 52880 60024 52886 60036
rect 567194 60024 567200 60036
rect 52880 59996 567200 60024
rect 52880 59984 52886 59996
rect 567194 59984 567200 59996
rect 567252 59984 567258 60036
rect 47578 59916 47584 59968
rect 47636 59956 47642 59968
rect 173894 59956 173900 59968
rect 47636 59928 173900 59956
rect 47636 59916 47642 59928
rect 173894 59916 173900 59928
rect 173952 59916 173958 59968
rect 202782 59916 202788 59968
rect 202840 59956 202846 59968
rect 446398 59956 446404 59968
rect 202840 59928 446404 59956
rect 202840 59916 202846 59928
rect 446398 59916 446404 59928
rect 446456 59916 446462 59968
rect 55950 59848 55956 59900
rect 56008 59888 56014 59900
rect 127158 59888 127164 59900
rect 56008 59860 127164 59888
rect 56008 59848 56014 59860
rect 127158 59848 127164 59860
rect 127216 59848 127222 59900
rect 168374 59888 168380 59900
rect 168335 59860 168380 59888
rect 168374 59848 168380 59860
rect 168432 59848 168438 59900
rect 211062 59888 211068 59900
rect 211023 59860 211068 59888
rect 211062 59848 211068 59860
rect 211120 59848 211126 59900
rect 218054 59888 218060 59900
rect 218015 59860 218060 59888
rect 218054 59848 218060 59860
rect 218112 59848 218118 59900
rect 224678 59888 224684 59900
rect 224639 59860 224684 59888
rect 224678 59848 224684 59860
rect 224736 59848 224742 59900
rect 227622 59848 227628 59900
rect 227680 59888 227686 59900
rect 442994 59888 443000 59900
rect 227680 59860 443000 59888
rect 227680 59848 227686 59860
rect 442994 59848 443000 59860
rect 443052 59848 443058 59900
rect 54846 59780 54852 59832
rect 54904 59820 54910 59832
rect 229186 59820 229192 59832
rect 54904 59792 229192 59820
rect 54904 59780 54910 59792
rect 229186 59780 229192 59792
rect 229244 59780 229250 59832
rect 235994 59820 236000 59832
rect 235955 59792 236000 59820
rect 235994 59780 236000 59792
rect 236052 59780 236058 59832
rect 248322 59780 248328 59832
rect 248380 59820 248386 59832
rect 441338 59820 441344 59832
rect 248380 59792 441344 59820
rect 248380 59780 248386 59792
rect 441338 59780 441344 59792
rect 441396 59780 441402 59832
rect 254026 59752 254032 59764
rect 253987 59724 254032 59752
rect 254026 59712 254032 59724
rect 254084 59712 254090 59764
rect 257982 59752 257988 59764
rect 257943 59724 257988 59752
rect 257982 59712 257988 59724
rect 258040 59712 258046 59764
rect 258074 59712 258080 59764
rect 258132 59752 258138 59764
rect 286962 59752 286968 59764
rect 258132 59724 258177 59752
rect 286923 59724 286968 59752
rect 258132 59712 258138 59724
rect 286962 59712 286968 59724
rect 287020 59712 287026 59764
rect 291102 59752 291108 59764
rect 291063 59724 291108 59752
rect 291102 59712 291108 59724
rect 291160 59712 291166 59764
rect 302234 59752 302240 59764
rect 302195 59724 302240 59752
rect 302234 59712 302240 59724
rect 302292 59712 302298 59764
rect 315942 59752 315948 59764
rect 315903 59724 315948 59752
rect 315942 59712 315948 59724
rect 316000 59712 316006 59764
rect 358814 59752 358820 59764
rect 358775 59724 358820 59752
rect 358814 59712 358820 59724
rect 358872 59712 358878 59764
rect 375374 59752 375380 59764
rect 375335 59724 375380 59752
rect 375374 59712 375380 59724
rect 375432 59712 375438 59764
rect 378042 59752 378048 59764
rect 378003 59724 378048 59752
rect 378042 59712 378048 59724
rect 378100 59712 378106 59764
rect 400122 59752 400128 59764
rect 400083 59724 400128 59752
rect 400122 59712 400128 59724
rect 400180 59712 400186 59764
rect 404262 59752 404268 59764
rect 404223 59724 404268 59752
rect 404262 59712 404268 59724
rect 404320 59712 404326 59764
rect 420914 59712 420920 59764
rect 420972 59752 420978 59764
rect 448606 59752 448612 59764
rect 420972 59724 448612 59752
rect 420972 59712 420978 59724
rect 448606 59712 448612 59724
rect 448664 59712 448670 59764
rect 375282 59684 375288 59696
rect 375243 59656 375288 59684
rect 375282 59644 375288 59656
rect 375340 59644 375346 59696
rect 414014 59644 414020 59696
rect 414072 59684 414078 59696
rect 439590 59684 439596 59696
rect 414072 59656 439596 59684
rect 414072 59644 414078 59656
rect 439590 59644 439596 59656
rect 439648 59644 439654 59696
rect 431862 59616 431868 59628
rect 431823 59588 431868 59616
rect 431862 59576 431868 59588
rect 431920 59576 431926 59628
rect 108942 59372 108948 59424
rect 109000 59412 109006 59424
rect 580166 59412 580172 59424
rect 109000 59384 580172 59412
rect 109000 59372 109006 59384
rect 580166 59372 580172 59384
rect 580224 59372 580230 59424
rect 2958 59304 2964 59356
rect 3016 59344 3022 59356
rect 25498 59344 25504 59356
rect 3016 59316 25504 59344
rect 3016 59304 3022 59316
rect 25498 59304 25504 59316
rect 25556 59304 25562 59356
rect 84470 59304 84476 59356
rect 84528 59344 84534 59356
rect 580442 59344 580448 59356
rect 84528 59316 580448 59344
rect 84528 59304 84534 59316
rect 580442 59304 580448 59316
rect 580500 59304 580506 59356
rect 114738 59236 114744 59288
rect 114796 59276 114802 59288
rect 580258 59276 580264 59288
rect 114796 59248 580264 59276
rect 114796 59236 114802 59248
rect 580258 59236 580264 59248
rect 580316 59236 580322 59288
rect 4890 59168 4896 59220
rect 4948 59208 4954 59220
rect 439314 59208 439320 59220
rect 4948 59180 439320 59208
rect 4948 59168 4954 59180
rect 439314 59168 439320 59180
rect 439372 59168 439378 59220
rect 3786 59100 3792 59152
rect 3844 59140 3850 59152
rect 320818 59140 320824 59152
rect 3844 59112 320824 59140
rect 3844 59100 3850 59112
rect 320818 59100 320824 59112
rect 320876 59100 320882 59152
rect 342714 59100 342720 59152
rect 342772 59140 342778 59152
rect 580626 59140 580632 59152
rect 342772 59112 580632 59140
rect 342772 59100 342778 59112
rect 580626 59100 580632 59112
rect 580684 59100 580690 59152
rect 3602 59032 3608 59084
rect 3660 59072 3666 59084
rect 238386 59072 238392 59084
rect 3660 59044 238392 59072
rect 3660 59032 3666 59044
rect 238386 59032 238392 59044
rect 238444 59032 238450 59084
rect 271230 59032 271236 59084
rect 271288 59072 271294 59084
rect 580810 59072 580816 59084
rect 271288 59044 580816 59072
rect 271288 59032 271294 59044
rect 580810 59032 580816 59044
rect 580868 59032 580874 59084
rect 24762 58964 24768 59016
rect 24820 59004 24826 59016
rect 293126 59004 293132 59016
rect 24820 58976 293132 59004
rect 24820 58964 24826 58976
rect 293126 58964 293132 58976
rect 293184 58964 293190 59016
rect 370406 58964 370412 59016
rect 370464 59004 370470 59016
rect 580350 59004 580356 59016
rect 370464 58976 580356 59004
rect 370464 58964 370470 58976
rect 580350 58964 580356 58976
rect 580408 58964 580414 59016
rect 171042 58896 171048 58948
rect 171100 58936 171106 58948
rect 446122 58936 446128 58948
rect 171100 58908 446128 58936
rect 171100 58896 171106 58908
rect 446122 58896 446128 58908
rect 446180 58896 446186 58948
rect 51258 58828 51264 58880
rect 51316 58868 51322 58880
rect 372614 58868 372620 58880
rect 51316 58840 372620 58868
rect 51316 58828 51322 58840
rect 372614 58828 372620 58840
rect 372672 58828 372678 58880
rect 402882 58828 402888 58880
rect 402940 58868 402946 58880
rect 440694 58868 440700 58880
rect 402940 58840 440700 58868
rect 402940 58828 402946 58840
rect 440694 58828 440700 58840
rect 440752 58828 440758 58880
rect 77202 58760 77208 58812
rect 77260 58800 77266 58812
rect 448054 58800 448060 58812
rect 77260 58772 448060 58800
rect 77260 58760 77266 58772
rect 448054 58760 448060 58772
rect 448112 58760 448118 58812
rect 52730 58692 52736 58744
rect 52788 58732 52794 58744
rect 524414 58732 524420 58744
rect 52788 58704 524420 58732
rect 52788 58692 52794 58704
rect 524414 58692 524420 58704
rect 524472 58692 524478 58744
rect 59078 58624 59084 58676
rect 59136 58664 59142 58676
rect 564526 58664 564532 58676
rect 59136 58636 564532 58664
rect 59136 58624 59142 58636
rect 564526 58624 564532 58636
rect 564584 58624 564590 58676
rect 188982 58556 188988 58608
rect 189040 58596 189046 58608
rect 446490 58596 446496 58608
rect 189040 58568 446496 58596
rect 189040 58556 189046 58568
rect 446490 58556 446496 58568
rect 446548 58556 446554 58608
rect 59722 58488 59728 58540
rect 59780 58528 59786 58540
rect 296714 58528 296720 58540
rect 59780 58500 296720 58528
rect 59780 58488 59786 58500
rect 296714 58488 296720 58500
rect 296772 58488 296778 58540
rect 345934 58488 345940 58540
rect 345992 58528 345998 58540
rect 462314 58528 462320 58540
rect 345992 58500 462320 58528
rect 345992 58488 345998 58500
rect 462314 58488 462320 58500
rect 462372 58488 462378 58540
rect 54202 58420 54208 58472
rect 54260 58460 54266 58472
rect 201494 58460 201500 58472
rect 54260 58432 201500 58460
rect 54260 58420 54266 58432
rect 201494 58420 201500 58432
rect 201552 58420 201558 58472
rect 233142 58420 233148 58472
rect 233200 58460 233206 58472
rect 439406 58460 439412 58472
rect 233200 58432 439412 58460
rect 233200 58420 233206 58432
rect 439406 58420 439412 58432
rect 439464 58420 439470 58472
rect 3878 58352 3884 58404
rect 3936 58392 3942 58404
rect 186222 58392 186228 58404
rect 3936 58364 186228 58392
rect 3936 58352 3942 58364
rect 186222 58352 186228 58364
rect 186280 58352 186286 58404
rect 422294 58352 422300 58404
rect 422352 58392 422358 58404
rect 450078 58392 450084 58404
rect 422352 58364 450084 58392
rect 422352 58352 422358 58364
rect 450078 58352 450084 58364
rect 450136 58352 450142 58404
rect 3510 58284 3516 58336
rect 3568 58324 3574 58336
rect 191374 58324 191380 58336
rect 3568 58296 191380 58324
rect 3568 58284 3574 58296
rect 191374 58284 191380 58296
rect 191432 58284 191438 58336
rect 434714 58284 434720 58336
rect 434772 58324 434778 58336
rect 452654 58324 452660 58336
rect 434772 58296 452660 58324
rect 434772 58284 434778 58296
rect 452654 58284 452660 58296
rect 452712 58284 452718 58336
rect 3418 57876 3424 57928
rect 3476 57916 3482 57928
rect 158530 57916 158536 57928
rect 3476 57888 158536 57916
rect 3476 57876 3482 57888
rect 158530 57876 158536 57888
rect 158588 57876 158594 57928
rect 172698 57876 172704 57928
rect 172756 57916 172762 57928
rect 173802 57916 173808 57928
rect 172756 57888 173808 57916
rect 172756 57876 172762 57888
rect 173802 57876 173808 57888
rect 173860 57876 173866 57928
rect 180426 57876 180432 57928
rect 180484 57916 180490 57928
rect 184934 57916 184940 57928
rect 180484 57888 184940 57916
rect 180484 57876 180490 57888
rect 184934 57876 184940 57888
rect 184992 57876 184998 57928
rect 188798 57876 188804 57928
rect 188856 57916 188862 57928
rect 307754 57916 307760 57928
rect 188856 57888 307760 57916
rect 188856 57876 188862 57888
rect 307754 57876 307760 57888
rect 307812 57876 307818 57928
rect 362862 57876 362868 57928
rect 362920 57916 362926 57928
rect 433518 57916 433524 57928
rect 362920 57888 433524 57916
rect 362920 57876 362926 57888
rect 433518 57876 433524 57888
rect 433576 57876 433582 57928
rect 73522 57808 73528 57860
rect 73580 57848 73586 57860
rect 74442 57848 74448 57860
rect 73580 57820 74448 57848
rect 73580 57808 73586 57820
rect 74442 57808 74448 57820
rect 74500 57808 74506 57860
rect 92842 57808 92848 57860
rect 92900 57848 92906 57860
rect 102226 57848 102232 57860
rect 92900 57820 102232 57848
rect 92900 57808 92906 57820
rect 102226 57808 102232 57820
rect 102284 57808 102290 57860
rect 123110 57808 123116 57860
rect 123168 57848 123174 57860
rect 226518 57848 226524 57860
rect 123168 57820 226524 57848
rect 123168 57808 123174 57820
rect 226518 57808 226524 57820
rect 226576 57808 226582 57860
rect 234522 57808 234528 57860
rect 234580 57848 234586 57860
rect 255130 57848 255136 57860
rect 234580 57820 255136 57848
rect 234580 57808 234586 57820
rect 255130 57808 255136 57820
rect 255188 57808 255194 57860
rect 279513 57851 279571 57857
rect 279513 57817 279525 57851
rect 279559 57848 279571 57851
rect 282178 57848 282184 57860
rect 279559 57820 282184 57848
rect 279559 57817 279571 57820
rect 279513 57811 279571 57817
rect 282178 57808 282184 57820
rect 282236 57808 282242 57860
rect 284202 57808 284208 57860
rect 284260 57848 284266 57860
rect 411622 57848 411628 57860
rect 284260 57820 411628 57848
rect 284260 57808 284266 57820
rect 411622 57808 411628 57820
rect 411680 57808 411686 57860
rect 419534 57808 419540 57860
rect 419592 57848 419598 57860
rect 444374 57848 444380 57860
rect 419592 57820 444380 57848
rect 419592 57808 419598 57820
rect 444374 57808 444380 57820
rect 444432 57808 444438 57860
rect 59998 57740 60004 57792
rect 60056 57780 60062 57792
rect 60056 57752 69704 57780
rect 60056 57740 60062 57752
rect 62574 57672 62580 57724
rect 62632 57712 62638 57724
rect 63310 57712 63316 57724
rect 62632 57684 63316 57712
rect 62632 57672 62638 57684
rect 63310 57672 63316 57684
rect 63368 57672 63374 57724
rect 67726 57672 67732 57724
rect 67784 57712 67790 57724
rect 68922 57712 68928 57724
rect 67784 57684 68928 57712
rect 67784 57672 67790 57684
rect 68922 57672 68928 57684
rect 68980 57672 68986 57724
rect 69676 57712 69704 57752
rect 69750 57740 69756 57792
rect 69808 57780 69814 57792
rect 101214 57780 101220 57792
rect 69808 57752 101220 57780
rect 69808 57740 69814 57752
rect 101214 57740 101220 57752
rect 101272 57740 101278 57792
rect 104802 57740 104808 57792
rect 104860 57780 104866 57792
rect 106366 57780 106372 57792
rect 104860 57752 106372 57780
rect 104860 57740 104866 57752
rect 106366 57740 106372 57752
rect 106424 57740 106430 57792
rect 112162 57740 112168 57792
rect 112220 57780 112226 57792
rect 112990 57780 112996 57792
rect 112220 57752 112996 57780
rect 112220 57740 112226 57752
rect 112990 57740 112996 57752
rect 113048 57740 113054 57792
rect 125505 57783 125563 57789
rect 125505 57780 125517 57783
rect 122806 57752 125517 57780
rect 81526 57712 81532 57724
rect 69676 57684 81532 57712
rect 81526 57672 81532 57684
rect 81584 57672 81590 57724
rect 87046 57672 87052 57724
rect 87104 57712 87110 57724
rect 122806 57712 122834 57752
rect 125505 57749 125517 57752
rect 125551 57749 125563 57783
rect 131482 57780 131488 57792
rect 125505 57743 125563 57749
rect 125704 57752 131488 57780
rect 87104 57684 122834 57712
rect 87104 57672 87110 57684
rect 28902 57604 28908 57656
rect 28960 57644 28966 57656
rect 125704 57644 125732 57752
rect 131482 57740 131488 57752
rect 131540 57740 131546 57792
rect 136634 57740 136640 57792
rect 136692 57780 136698 57792
rect 136692 57752 140176 57780
rect 136692 57740 136698 57752
rect 125781 57715 125839 57721
rect 125781 57681 125793 57715
rect 125827 57712 125839 57715
rect 139949 57715 140007 57721
rect 139949 57712 139961 57715
rect 125827 57684 139961 57712
rect 125827 57681 125839 57684
rect 125781 57675 125839 57681
rect 139949 57681 139961 57684
rect 139995 57681 140007 57715
rect 139949 57675 140007 57681
rect 28960 57616 125732 57644
rect 28960 57604 28966 57616
rect 139210 57604 139216 57656
rect 139268 57644 139274 57656
rect 140038 57644 140044 57656
rect 139268 57616 140044 57644
rect 139268 57604 139274 57616
rect 140038 57604 140044 57616
rect 140096 57604 140102 57656
rect 140148 57644 140176 57752
rect 142430 57740 142436 57792
rect 142488 57780 142494 57792
rect 143442 57780 143448 57792
rect 142488 57752 143448 57780
rect 142488 57740 142494 57752
rect 143442 57740 143448 57752
rect 143500 57740 143506 57792
rect 145006 57740 145012 57792
rect 145064 57780 145070 57792
rect 146202 57780 146208 57792
rect 145064 57752 146208 57780
rect 145064 57740 145070 57752
rect 146202 57740 146208 57752
rect 146260 57740 146266 57792
rect 148962 57740 148968 57792
rect 149020 57780 149026 57792
rect 287974 57780 287980 57792
rect 149020 57752 287980 57780
rect 149020 57740 149026 57752
rect 287974 57740 287980 57752
rect 288032 57740 288038 57792
rect 326614 57740 326620 57792
rect 326672 57780 326678 57792
rect 439038 57780 439044 57792
rect 326672 57752 439044 57780
rect 326672 57740 326678 57752
rect 439038 57740 439044 57752
rect 439096 57740 439102 57792
rect 140225 57715 140283 57721
rect 140225 57681 140237 57715
rect 140271 57712 140283 57715
rect 191834 57712 191840 57724
rect 140271 57684 191840 57712
rect 140271 57681 140283 57684
rect 140225 57675 140283 57681
rect 191834 57672 191840 57684
rect 191892 57672 191898 57724
rect 194594 57672 194600 57724
rect 194652 57712 194658 57724
rect 195882 57712 195888 57724
rect 194652 57684 195888 57712
rect 194652 57672 194658 57684
rect 195882 57672 195888 57684
rect 195940 57672 195946 57724
rect 209866 57672 209872 57724
rect 209924 57712 209930 57724
rect 210694 57712 210700 57724
rect 209924 57684 210700 57712
rect 209924 57672 209930 57684
rect 210694 57672 210700 57684
rect 210752 57672 210758 57724
rect 213822 57672 213828 57724
rect 213880 57712 213886 57724
rect 353662 57712 353668 57724
rect 213880 57684 353668 57712
rect 213880 57672 213886 57684
rect 353662 57672 353668 57684
rect 353720 57672 353726 57724
rect 376202 57672 376208 57724
rect 376260 57712 376266 57724
rect 381538 57712 381544 57724
rect 376260 57684 381544 57712
rect 376260 57672 376266 57684
rect 381538 57672 381544 57684
rect 381596 57672 381602 57724
rect 387150 57672 387156 57724
rect 387208 57712 387214 57724
rect 463694 57712 463700 57724
rect 387208 57684 463700 57712
rect 387208 57672 387214 57684
rect 463694 57672 463700 57684
rect 463752 57672 463758 57724
rect 287054 57644 287060 57656
rect 140148 57616 287060 57644
rect 287054 57604 287060 57616
rect 287112 57604 287118 57656
rect 323394 57604 323400 57656
rect 323452 57644 323458 57656
rect 324222 57644 324228 57656
rect 323452 57616 324228 57644
rect 323452 57604 323458 57616
rect 324222 57604 324228 57616
rect 324280 57604 324286 57656
rect 343542 57604 343548 57656
rect 343600 57644 343606 57656
rect 389726 57644 389732 57656
rect 343600 57616 389732 57644
rect 343600 57604 343606 57616
rect 389726 57604 389732 57616
rect 389784 57604 389790 57656
rect 403250 57604 403256 57656
rect 403308 57644 403314 57656
rect 407758 57644 407764 57656
rect 403308 57616 407764 57644
rect 403308 57604 403314 57616
rect 407758 57604 407764 57616
rect 407816 57604 407822 57656
rect 409509 57647 409567 57653
rect 409509 57613 409521 57647
rect 409555 57644 409567 57647
rect 542998 57644 543004 57656
rect 409555 57616 543004 57644
rect 409555 57613 409567 57616
rect 409509 57607 409567 57613
rect 542998 57604 543004 57616
rect 543056 57604 543062 57656
rect 13722 57536 13728 57588
rect 13780 57576 13786 57588
rect 127894 57576 127900 57588
rect 13780 57548 127900 57576
rect 13780 57536 13786 57548
rect 127894 57536 127900 57548
rect 127952 57536 127958 57588
rect 128262 57536 128268 57588
rect 128320 57576 128326 57588
rect 279513 57579 279571 57585
rect 279513 57576 279525 57579
rect 128320 57548 279525 57576
rect 128320 57536 128326 57548
rect 279513 57545 279525 57548
rect 279559 57545 279571 57579
rect 279513 57539 279571 57545
rect 279602 57536 279608 57588
rect 279660 57576 279666 57588
rect 282178 57576 282184 57588
rect 279660 57548 282184 57576
rect 279660 57536 279666 57548
rect 282178 57536 282184 57548
rect 282236 57536 282242 57588
rect 356882 57536 356888 57588
rect 356940 57576 356946 57588
rect 364334 57576 364340 57588
rect 356940 57548 364340 57576
rect 356940 57536 356946 57548
rect 364334 57536 364340 57548
rect 364392 57536 364398 57588
rect 367830 57536 367836 57588
rect 367888 57576 367894 57588
rect 518250 57576 518256 57588
rect 367888 57548 518256 57576
rect 367888 57536 367894 57548
rect 518250 57536 518256 57548
rect 518308 57536 518314 57588
rect 34422 57468 34428 57520
rect 34480 57508 34486 57520
rect 202966 57508 202972 57520
rect 34480 57480 202972 57508
rect 34480 57468 34486 57480
rect 202966 57468 202972 57480
rect 203024 57468 203030 57520
rect 233234 57468 233240 57520
rect 233292 57508 233298 57520
rect 234430 57508 234436 57520
rect 233292 57480 234436 57508
rect 233292 57468 233298 57480
rect 234430 57468 234436 57480
rect 234488 57468 234494 57520
rect 240962 57468 240968 57520
rect 241020 57508 241026 57520
rect 298738 57508 298744 57520
rect 241020 57480 298744 57508
rect 241020 57468 241026 57480
rect 298738 57468 298744 57480
rect 298796 57468 298802 57520
rect 309870 57468 309876 57520
rect 309928 57508 309934 57520
rect 320818 57508 320824 57520
rect 309928 57480 320824 57508
rect 309928 57468 309934 57480
rect 320818 57468 320824 57480
rect 320876 57468 320882 57520
rect 329190 57468 329196 57520
rect 329248 57508 329254 57520
rect 531958 57508 531964 57520
rect 329248 57480 531964 57508
rect 329248 57468 329254 57480
rect 531958 57468 531964 57480
rect 532016 57468 532022 57520
rect 55030 57400 55036 57452
rect 55088 57440 55094 57452
rect 244274 57440 244280 57452
rect 55088 57412 244280 57440
rect 55088 57400 55094 57412
rect 244274 57400 244280 57412
rect 244332 57400 244338 57452
rect 273162 57400 273168 57452
rect 273220 57440 273226 57452
rect 296346 57440 296352 57452
rect 273220 57412 296352 57440
rect 273220 57400 273226 57412
rect 296346 57400 296352 57412
rect 296404 57400 296410 57452
rect 301498 57400 301504 57452
rect 301556 57440 301562 57452
rect 509878 57440 509884 57452
rect 301556 57412 509884 57440
rect 301556 57400 301562 57412
rect 509878 57400 509884 57412
rect 509936 57400 509942 57452
rect 37182 57332 37188 57384
rect 37240 57372 37246 57384
rect 81894 57372 81900 57384
rect 37240 57344 81900 57372
rect 37240 57332 37246 57344
rect 81894 57332 81900 57344
rect 81952 57332 81958 57384
rect 89622 57332 89628 57384
rect 89680 57372 89686 57384
rect 299474 57372 299480 57384
rect 89680 57344 299480 57372
rect 89680 57332 89686 57344
rect 299474 57332 299480 57344
rect 299532 57332 299538 57384
rect 304718 57332 304724 57384
rect 304776 57372 304782 57384
rect 523678 57372 523684 57384
rect 304776 57344 523684 57372
rect 304776 57332 304782 57344
rect 523678 57332 523684 57344
rect 523736 57332 523742 57384
rect 10962 57264 10968 57316
rect 11020 57304 11026 57316
rect 95418 57304 95424 57316
rect 11020 57276 95424 57304
rect 11020 57264 11026 57276
rect 95418 57264 95424 57276
rect 95476 57264 95482 57316
rect 119890 57264 119896 57316
rect 119948 57304 119954 57316
rect 447778 57304 447784 57316
rect 119948 57276 447784 57304
rect 119948 57264 119954 57276
rect 447778 57264 447784 57276
rect 447836 57264 447842 57316
rect 22002 57196 22008 57248
rect 22060 57236 22066 57248
rect 404449 57239 404507 57245
rect 404449 57236 404461 57239
rect 22060 57208 404461 57236
rect 22060 57196 22066 57208
rect 404449 57205 404461 57208
rect 404495 57205 404507 57239
rect 404449 57199 404507 57205
rect 406470 57196 406476 57248
rect 406528 57236 406534 57248
rect 409509 57239 409567 57245
rect 409509 57236 409521 57239
rect 406528 57208 409521 57236
rect 406528 57196 406534 57208
rect 409509 57205 409521 57208
rect 409555 57205 409567 57239
rect 409509 57199 409567 57205
rect 414198 57196 414204 57248
rect 414256 57236 414262 57248
rect 448606 57236 448612 57248
rect 414256 57208 448612 57236
rect 414256 57196 414262 57208
rect 448606 57196 448612 57208
rect 448664 57196 448670 57248
rect 63402 57128 63408 57180
rect 63460 57168 63466 57180
rect 155954 57168 155960 57180
rect 63460 57140 155960 57168
rect 63460 57128 63466 57140
rect 155954 57128 155960 57140
rect 156012 57128 156018 57180
rect 175274 57128 175280 57180
rect 175332 57168 175338 57180
rect 291194 57168 291200 57180
rect 175332 57140 291200 57168
rect 175332 57128 175338 57140
rect 291194 57128 291200 57140
rect 291252 57128 291258 57180
rect 393222 57128 393228 57180
rect 393280 57168 393286 57180
rect 449250 57168 449256 57180
rect 393280 57140 449256 57168
rect 393280 57128 393286 57140
rect 449250 57128 449256 57140
rect 449308 57128 449314 57180
rect 103790 57060 103796 57112
rect 103848 57100 103854 57112
rect 205634 57100 205640 57112
rect 103848 57072 205640 57100
rect 103848 57060 103854 57072
rect 205634 57060 205640 57072
rect 205692 57060 205698 57112
rect 220722 57060 220728 57112
rect 220780 57100 220786 57112
rect 331766 57100 331772 57112
rect 220780 57072 331772 57100
rect 220780 57060 220786 57072
rect 331766 57060 331772 57072
rect 331824 57060 331830 57112
rect 407022 57060 407028 57112
rect 407080 57100 407086 57112
rect 441062 57100 441068 57112
rect 407080 57072 441068 57100
rect 407080 57060 407086 57072
rect 441062 57060 441068 57072
rect 441120 57060 441126 57112
rect 100662 56992 100668 57044
rect 100720 57032 100726 57044
rect 150158 57032 150164 57044
rect 100720 57004 150164 57032
rect 100720 56992 100726 57004
rect 150158 56992 150164 57004
rect 150216 56992 150222 57044
rect 182082 56992 182088 57044
rect 182140 57032 182146 57044
rect 285398 57032 285404 57044
rect 182140 57004 285404 57032
rect 182140 56992 182146 57004
rect 285398 56992 285404 57004
rect 285456 56992 285462 57044
rect 400674 56992 400680 57044
rect 400732 57032 400738 57044
rect 416774 57032 416780 57044
rect 400732 57004 416780 57032
rect 400732 56992 400738 57004
rect 416774 56992 416780 57004
rect 416832 56992 416838 57044
rect 419994 56992 420000 57044
rect 420052 57032 420058 57044
rect 429194 57032 429200 57044
rect 420052 57004 429200 57032
rect 420052 56992 420058 57004
rect 429194 56992 429200 57004
rect 429252 56992 429258 57044
rect 125686 56924 125692 56976
rect 125744 56964 125750 56976
rect 126882 56964 126888 56976
rect 125744 56936 126888 56964
rect 125744 56924 125750 56936
rect 126882 56924 126888 56936
rect 126940 56924 126946 56976
rect 134058 56924 134064 56976
rect 134116 56964 134122 56976
rect 157334 56964 157340 56976
rect 134116 56936 157340 56964
rect 134116 56924 134122 56936
rect 157334 56924 157340 56936
rect 157392 56924 157398 56976
rect 160002 56924 160008 56976
rect 160060 56964 160066 56976
rect 249334 56964 249340 56976
rect 160060 56936 249340 56964
rect 160060 56924 160066 56936
rect 249334 56924 249340 56936
rect 249392 56924 249398 56976
rect 404449 56967 404507 56973
rect 404449 56933 404461 56967
rect 404495 56964 404507 56967
rect 409046 56964 409052 56976
rect 404495 56936 409052 56964
rect 404495 56933 404507 56936
rect 404449 56927 404507 56933
rect 409046 56924 409052 56936
rect 409104 56924 409110 56976
rect 76098 56856 76104 56908
rect 76156 56896 76162 56908
rect 83458 56896 83464 56908
rect 76156 56868 83464 56896
rect 76156 56856 76162 56868
rect 83458 56856 83464 56868
rect 83516 56856 83522 56908
rect 113082 56856 113088 56908
rect 113140 56896 113146 56908
rect 197170 56896 197176 56908
rect 113140 56868 197176 56896
rect 113140 56856 113146 56868
rect 197170 56856 197176 56868
rect 197228 56856 197234 56908
rect 212442 56856 212448 56908
rect 212500 56896 212506 56908
rect 251910 56896 251916 56908
rect 212500 56868 251916 56896
rect 212500 56856 212506 56868
rect 251910 56856 251916 56868
rect 251968 56856 251974 56908
rect 164142 56788 164148 56840
rect 164200 56828 164206 56840
rect 230014 56828 230020 56840
rect 164200 56800 230020 56828
rect 164200 56788 164206 56800
rect 230014 56788 230020 56800
rect 230072 56788 230078 56840
rect 97994 56720 98000 56772
rect 98052 56760 98058 56772
rect 99190 56760 99196 56772
rect 98052 56732 99196 56760
rect 98052 56720 98058 56732
rect 99190 56720 99196 56732
rect 99248 56720 99254 56772
rect 129642 56720 129648 56772
rect 129700 56760 129706 56772
rect 164326 56760 164332 56772
rect 129700 56732 164332 56760
rect 129700 56720 129706 56732
rect 164326 56720 164332 56732
rect 164384 56720 164390 56772
rect 183646 56720 183652 56772
rect 183704 56760 183710 56772
rect 194686 56760 194692 56772
rect 183704 56732 194692 56760
rect 183704 56720 183710 56732
rect 194686 56720 194692 56732
rect 194744 56720 194750 56772
rect 65150 56652 65156 56704
rect 65208 56692 65214 56704
rect 66070 56692 66076 56704
rect 65208 56664 66076 56692
rect 65208 56652 65214 56664
rect 66070 56652 66076 56664
rect 66128 56652 66134 56704
rect 117314 56584 117320 56636
rect 117372 56624 117378 56636
rect 123478 56624 123484 56636
rect 117372 56596 123484 56624
rect 117372 56584 117378 56596
rect 123478 56584 123484 56596
rect 123536 56584 123542 56636
rect 295978 56584 295984 56636
rect 296036 56624 296042 56636
rect 298922 56624 298928 56636
rect 296036 56596 298928 56624
rect 296036 56584 296042 56596
rect 298922 56584 298928 56596
rect 298980 56584 298986 56636
rect 353202 56516 353208 56568
rect 353260 56556 353266 56568
rect 451274 56556 451280 56568
rect 353260 56528 451280 56556
rect 353260 56516 353266 56528
rect 451274 56516 451280 56528
rect 451332 56516 451338 56568
rect 58158 56448 58164 56500
rect 58216 56488 58222 56500
rect 200114 56488 200120 56500
rect 58216 56460 200120 56488
rect 58216 56448 58222 56460
rect 200114 56448 200120 56460
rect 200172 56448 200178 56500
rect 274542 56448 274548 56500
rect 274600 56488 274606 56500
rect 441430 56488 441436 56500
rect 274600 56460 441436 56488
rect 274600 56448 274606 56460
rect 441430 56448 441436 56460
rect 441488 56448 441494 56500
rect 49234 56380 49240 56432
rect 49292 56420 49298 56432
rect 178034 56420 178040 56432
rect 49292 56392 178040 56420
rect 49292 56380 49298 56392
rect 178034 56380 178040 56392
rect 178092 56380 178098 56432
rect 191742 56380 191748 56432
rect 191800 56420 191806 56432
rect 450630 56420 450636 56432
rect 191800 56392 450636 56420
rect 191800 56380 191806 56392
rect 450630 56380 450636 56392
rect 450688 56380 450694 56432
rect 58250 56312 58256 56364
rect 58308 56352 58314 56364
rect 324314 56352 324320 56364
rect 58308 56324 324320 56352
rect 58308 56312 58314 56324
rect 324314 56312 324320 56324
rect 324372 56312 324378 56364
rect 346302 56312 346308 56364
rect 346360 56352 346366 56364
rect 450446 56352 450452 56364
rect 346360 56324 450452 56352
rect 346360 56312 346366 56324
rect 450446 56312 450452 56324
rect 450504 56312 450510 56364
rect 59814 56244 59820 56296
rect 59872 56284 59878 56296
rect 423674 56284 423680 56296
rect 59872 56256 423680 56284
rect 59872 56244 59878 56256
rect 423674 56244 423680 56256
rect 423732 56244 423738 56296
rect 433242 56244 433248 56296
rect 433300 56284 433306 56296
rect 454218 56284 454224 56296
rect 433300 56256 454224 56284
rect 433300 56244 433306 56256
rect 454218 56244 454224 56256
rect 454276 56244 454282 56296
rect 66162 56176 66168 56228
rect 66220 56216 66226 56228
rect 447594 56216 447600 56228
rect 66220 56188 447600 56216
rect 66220 56176 66226 56188
rect 447594 56176 447600 56188
rect 447652 56176 447658 56228
rect 56962 56108 56968 56160
rect 57020 56148 57026 56160
rect 472710 56148 472716 56160
rect 57020 56120 472716 56148
rect 57020 56108 57026 56120
rect 472710 56108 472716 56120
rect 472768 56108 472774 56160
rect 3418 56040 3424 56092
rect 3476 56080 3482 56092
rect 440050 56080 440056 56092
rect 3476 56052 440056 56080
rect 3476 56040 3482 56052
rect 440050 56040 440056 56052
rect 440108 56040 440114 56092
rect 50154 55972 50160 56024
rect 50212 56012 50218 56024
rect 527174 56012 527180 56024
rect 50212 55984 527180 56012
rect 50212 55972 50218 55984
rect 527174 55972 527180 55984
rect 527232 55972 527238 56024
rect 49510 55904 49516 55956
rect 49568 55944 49574 55956
rect 568574 55944 568580 55956
rect 49568 55916 568580 55944
rect 49568 55904 49574 55916
rect 568574 55904 568580 55916
rect 568632 55904 568638 55956
rect 45462 55836 45468 55888
rect 45520 55876 45526 55888
rect 580258 55876 580264 55888
rect 45520 55848 580264 55876
rect 45520 55836 45526 55848
rect 580258 55836 580264 55848
rect 580316 55836 580322 55888
rect 397362 55768 397368 55820
rect 397420 55808 397426 55820
rect 445110 55808 445116 55820
rect 397420 55780 445116 55808
rect 397420 55768 397426 55780
rect 445110 55768 445116 55780
rect 445168 55768 445174 55820
rect 429102 55700 429108 55752
rect 429160 55740 429166 55752
rect 446674 55740 446680 55752
rect 429160 55712 446680 55740
rect 429160 55700 429166 55712
rect 446674 55700 446680 55712
rect 446732 55700 446738 55752
rect 249702 55020 249708 55072
rect 249760 55060 249766 55072
rect 451550 55060 451556 55072
rect 249760 55032 451556 55060
rect 249760 55020 249766 55032
rect 451550 55020 451556 55032
rect 451608 55020 451614 55072
rect 49142 54952 49148 55004
rect 49200 54992 49206 55004
rect 255314 54992 255320 55004
rect 49200 54964 255320 54992
rect 49200 54952 49206 54964
rect 255314 54952 255320 54964
rect 255372 54952 255378 55004
rect 47946 54884 47952 54936
rect 48004 54924 48010 54936
rect 284294 54924 284300 54936
rect 48004 54896 284300 54924
rect 48004 54884 48010 54896
rect 284294 54884 284300 54896
rect 284352 54884 284358 54936
rect 400030 54884 400036 54936
rect 400088 54924 400094 54936
rect 444742 54924 444748 54936
rect 400088 54896 444748 54924
rect 400088 54884 400094 54896
rect 444742 54884 444748 54896
rect 444800 54884 444806 54936
rect 180702 54816 180708 54868
rect 180760 54856 180766 54868
rect 451366 54856 451372 54868
rect 180760 54828 451372 54856
rect 180760 54816 180766 54828
rect 451366 54816 451372 54828
rect 451424 54816 451430 54868
rect 59630 54748 59636 54800
rect 59688 54788 59694 54800
rect 349154 54788 349160 54800
rect 59688 54760 349160 54788
rect 59688 54748 59694 54760
rect 349154 54748 349160 54760
rect 349212 54748 349218 54800
rect 371142 54748 371148 54800
rect 371200 54788 371206 54800
rect 452930 54788 452936 54800
rect 371200 54760 452936 54788
rect 371200 54748 371206 54760
rect 452930 54748 452936 54760
rect 452988 54748 452994 54800
rect 135162 54680 135168 54732
rect 135220 54720 135226 54732
rect 439958 54720 439964 54732
rect 135220 54692 439964 54720
rect 135220 54680 135226 54692
rect 439958 54680 439964 54692
rect 440016 54680 440022 54732
rect 49326 54612 49332 54664
rect 49384 54652 49390 54664
rect 540974 54652 540980 54664
rect 49384 54624 540980 54652
rect 49384 54612 49390 54624
rect 540974 54612 540980 54624
rect 541032 54612 541038 54664
rect 46750 54544 46756 54596
rect 46808 54584 46814 54596
rect 557534 54584 557540 54596
rect 46808 54556 557540 54584
rect 46808 54544 46814 54556
rect 557534 54544 557540 54556
rect 557592 54544 557598 54596
rect 47762 54476 47768 54528
rect 47820 54516 47826 54528
rect 575474 54516 575480 54528
rect 47820 54488 575480 54516
rect 47820 54476 47826 54488
rect 575474 54476 575480 54488
rect 575532 54476 575538 54528
rect 295242 53524 295248 53576
rect 295300 53564 295306 53576
rect 445018 53564 445024 53576
rect 295300 53536 445024 53564
rect 295300 53524 295306 53536
rect 445018 53524 445024 53536
rect 445076 53524 445082 53576
rect 44910 53456 44916 53508
rect 44968 53496 44974 53508
rect 209774 53496 209780 53508
rect 44968 53468 209780 53496
rect 44968 53456 44974 53468
rect 209774 53456 209780 53468
rect 209832 53456 209838 53508
rect 285582 53456 285588 53508
rect 285640 53496 285646 53508
rect 446582 53496 446588 53508
rect 285640 53468 446588 53496
rect 285640 53456 285646 53468
rect 446582 53456 446588 53468
rect 446640 53456 446646 53508
rect 184842 53388 184848 53440
rect 184900 53428 184906 53440
rect 439774 53428 439780 53440
rect 184900 53400 439780 53428
rect 184900 53388 184906 53400
rect 439774 53388 439780 53400
rect 439832 53388 439838 53440
rect 43990 53320 43996 53372
rect 44048 53360 44054 53372
rect 338114 53360 338120 53372
rect 44048 53332 338120 53360
rect 44048 53320 44054 53332
rect 338114 53320 338120 53332
rect 338172 53320 338178 53372
rect 354582 53320 354588 53372
rect 354640 53360 354646 53372
rect 453114 53360 453120 53372
rect 354640 53332 453120 53360
rect 354640 53320 354646 53332
rect 453114 53320 453120 53332
rect 453172 53320 453178 53372
rect 51166 53252 51172 53304
rect 51224 53292 51230 53304
rect 365714 53292 365720 53304
rect 51224 53264 365720 53292
rect 51224 53252 51230 53264
rect 365714 53252 365720 53264
rect 365772 53252 365778 53304
rect 369762 53252 369768 53304
rect 369820 53292 369826 53304
rect 450538 53292 450544 53304
rect 369820 53264 450544 53292
rect 369820 53252 369826 53264
rect 450538 53252 450544 53264
rect 450596 53252 450602 53304
rect 46474 53184 46480 53236
rect 46532 53224 46538 53236
rect 386414 53224 386420 53236
rect 46532 53196 386420 53224
rect 46532 53184 46538 53196
rect 386414 53184 386420 53196
rect 386472 53184 386478 53236
rect 47486 53116 47492 53168
rect 47544 53156 47550 53168
rect 409874 53156 409880 53168
rect 47544 53128 409880 53156
rect 47544 53116 47550 53128
rect 409874 53116 409880 53128
rect 409932 53116 409938 53168
rect 52546 53048 52552 53100
rect 52604 53088 52610 53100
rect 470594 53088 470600 53100
rect 52604 53060 470600 53088
rect 52604 53048 52610 53060
rect 470594 53048 470600 53060
rect 470652 53048 470658 53100
rect 213914 52028 213920 52080
rect 213972 52068 213978 52080
rect 367094 52068 367100 52080
rect 213972 52040 367100 52068
rect 213972 52028 213978 52040
rect 367094 52028 367100 52040
rect 367152 52028 367158 52080
rect 43898 51960 43904 52012
rect 43956 52000 43962 52012
rect 288434 52000 288440 52012
rect 43956 51972 288440 52000
rect 43956 51960 43962 51972
rect 288434 51960 288440 51972
rect 288492 51960 288498 52012
rect 310422 51960 310428 52012
rect 310480 52000 310486 52012
rect 445846 52000 445852 52012
rect 310480 51972 445852 52000
rect 310480 51960 310486 51972
rect 445846 51960 445852 51972
rect 445904 51960 445910 52012
rect 132402 51892 132408 51944
rect 132460 51932 132466 51944
rect 451642 51932 451648 51944
rect 132460 51904 451648 51932
rect 132460 51892 132466 51904
rect 451642 51892 451648 51904
rect 451700 51892 451706 51944
rect 45094 51824 45100 51876
rect 45152 51864 45158 51876
rect 382274 51864 382280 51876
rect 45152 51836 382280 51864
rect 45152 51824 45158 51836
rect 382274 51824 382280 51836
rect 382332 51824 382338 51876
rect 209866 51756 209872 51808
rect 209924 51796 209930 51808
rect 555418 51796 555424 51808
rect 209924 51768 555424 51796
rect 209924 51756 209930 51768
rect 555418 51756 555424 51768
rect 555476 51756 555482 51808
rect 46290 51688 46296 51740
rect 46348 51728 46354 51740
rect 423766 51728 423772 51740
rect 46348 51700 423772 51728
rect 46348 51688 46354 51700
rect 423766 51688 423772 51700
rect 423824 51688 423830 51740
rect 111702 50532 111708 50584
rect 111760 50572 111766 50584
rect 457070 50572 457076 50584
rect 111760 50544 457076 50572
rect 111760 50532 111766 50544
rect 457070 50532 457076 50544
rect 457128 50532 457134 50584
rect 95142 50464 95148 50516
rect 95200 50504 95206 50516
rect 454402 50504 454408 50516
rect 95200 50476 454408 50504
rect 95200 50464 95206 50476
rect 454402 50464 454408 50476
rect 454460 50464 454466 50516
rect 62022 50396 62028 50448
rect 62080 50436 62086 50448
rect 447502 50436 447508 50448
rect 62080 50408 447508 50436
rect 62080 50396 62086 50408
rect 447502 50396 447508 50408
rect 447560 50396 447566 50448
rect 53374 50328 53380 50380
rect 53432 50368 53438 50380
rect 485774 50368 485780 50380
rect 53432 50340 485780 50368
rect 53432 50328 53438 50340
rect 485774 50328 485780 50340
rect 485832 50328 485838 50380
rect 79962 48968 79968 49020
rect 80020 49008 80026 49020
rect 446766 49008 446772 49020
rect 80020 48980 446772 49008
rect 80020 48968 80026 48980
rect 446766 48968 446772 48980
rect 446824 48968 446830 49020
rect 54938 47540 54944 47592
rect 54996 47580 55002 47592
rect 129734 47580 129740 47592
rect 54996 47552 129740 47580
rect 54996 47540 55002 47552
rect 129734 47540 129740 47552
rect 129792 47540 129798 47592
rect 166902 47540 166908 47592
rect 166960 47580 166966 47592
rect 492674 47580 492680 47592
rect 166960 47552 492680 47580
rect 166960 47540 166966 47552
rect 492674 47540 492680 47552
rect 492732 47540 492738 47592
rect 99190 46860 99196 46912
rect 99248 46900 99254 46912
rect 580166 46900 580172 46912
rect 99248 46872 580172 46900
rect 99248 46860 99254 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 245654 45540 245660 45552
rect 3568 45512 245660 45540
rect 3568 45500 3574 45512
rect 245654 45500 245660 45512
rect 245712 45500 245718 45552
rect 37090 39380 37096 39432
rect 37148 39420 37154 39432
rect 448790 39420 448796 39432
rect 37148 39392 448796 39420
rect 37148 39380 37154 39392
rect 448790 39380 448796 39392
rect 448848 39380 448854 39432
rect 56042 39312 56048 39364
rect 56100 39352 56106 39364
rect 476114 39352 476120 39364
rect 56100 39324 476120 39352
rect 56100 39312 56106 39324
rect 476114 39312 476120 39324
rect 476172 39312 476178 39364
rect 472618 33056 472624 33108
rect 472676 33096 472682 33108
rect 580166 33096 580172 33108
rect 472676 33068 580172 33096
rect 472676 33056 472682 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 58342 28228 58348 28280
rect 58400 28268 58406 28280
rect 220906 28268 220912 28280
rect 58400 28240 220912 28268
rect 58400 28228 58406 28240
rect 220906 28228 220912 28240
rect 220964 28228 220970 28280
rect 277302 28228 277308 28280
rect 277360 28268 277366 28280
rect 536098 28268 536104 28280
rect 277360 28240 536104 28268
rect 277360 28228 277366 28240
rect 536098 28228 536104 28240
rect 536156 28228 536162 28280
rect 299382 26868 299388 26920
rect 299440 26908 299446 26920
rect 453022 26908 453028 26920
rect 299440 26880 453028 26908
rect 299440 26868 299446 26880
rect 453022 26868 453028 26880
rect 453080 26868 453086 26920
rect 140038 25508 140044 25560
rect 140096 25548 140102 25560
rect 528554 25548 528560 25560
rect 140096 25520 528560 25548
rect 140096 25508 140102 25520
rect 528554 25508 528560 25520
rect 528612 25508 528618 25560
rect 209682 22788 209688 22840
rect 209740 22828 209746 22840
rect 454310 22828 454316 22840
rect 209740 22800 454316 22828
rect 209740 22788 209746 22800
rect 454310 22788 454316 22800
rect 454368 22788 454374 22840
rect 46382 22720 46388 22772
rect 46440 22760 46446 22772
rect 325694 22760 325700 22772
rect 46440 22732 325700 22760
rect 46440 22720 46446 22732
rect 325694 22720 325700 22732
rect 325752 22720 325758 22772
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 436094 20652 436100 20664
rect 3476 20624 436100 20652
rect 3476 20612 3482 20624
rect 436094 20612 436100 20624
rect 436152 20612 436158 20664
rect 282178 17212 282184 17264
rect 282236 17252 282242 17264
rect 328454 17252 328460 17264
rect 282236 17224 328460 17252
rect 282236 17212 282242 17224
rect 328454 17212 328460 17224
rect 328512 17212 328518 17264
rect 335262 17212 335268 17264
rect 335320 17252 335326 17264
rect 500218 17252 500224 17264
rect 335320 17224 500224 17252
rect 335320 17212 335326 17224
rect 500218 17212 500224 17224
rect 500276 17212 500282 17264
rect 45278 15988 45284 16040
rect 45336 16028 45342 16040
rect 214466 16028 214472 16040
rect 45336 16000 214472 16028
rect 45336 15988 45342 16000
rect 214466 15988 214472 16000
rect 214524 15988 214530 16040
rect 216582 15988 216588 16040
rect 216640 16028 216646 16040
rect 407206 16028 407212 16040
rect 216640 16000 407212 16028
rect 216640 15988 216646 16000
rect 407206 15988 407212 16000
rect 407264 15988 407270 16040
rect 173802 15920 173808 15972
rect 173860 15960 173866 15972
rect 382366 15960 382372 15972
rect 173860 15932 382372 15960
rect 173860 15920 173866 15932
rect 382366 15920 382372 15932
rect 382424 15920 382430 15972
rect 123478 15852 123484 15904
rect 123536 15892 123542 15904
rect 339862 15892 339868 15904
rect 123536 15864 339868 15892
rect 123536 15852 123542 15864
rect 339862 15852 339868 15864
rect 339920 15852 339926 15904
rect 384758 15852 384764 15904
rect 384816 15892 384822 15904
rect 439866 15892 439872 15904
rect 384816 15864 439872 15892
rect 384816 15852 384822 15864
rect 439866 15852 439872 15864
rect 439924 15852 439930 15904
rect 260742 14696 260748 14748
rect 260800 14736 260806 14748
rect 361114 14736 361120 14748
rect 260800 14708 361120 14736
rect 260800 14696 260806 14708
rect 361114 14696 361120 14708
rect 361172 14696 361178 14748
rect 269022 14628 269028 14680
rect 269080 14668 269086 14680
rect 389450 14668 389456 14680
rect 269080 14640 389456 14668
rect 269080 14628 269086 14640
rect 389450 14628 389456 14640
rect 389508 14628 389514 14680
rect 176562 14560 176568 14612
rect 176620 14600 176626 14612
rect 450170 14600 450176 14612
rect 176620 14572 450176 14600
rect 176620 14560 176626 14572
rect 450170 14560 450176 14572
rect 450228 14560 450234 14612
rect 43806 14492 43812 14544
rect 43864 14532 43870 14544
rect 379974 14532 379980 14544
rect 43864 14504 379980 14532
rect 43864 14492 43870 14504
rect 379974 14492 379980 14504
rect 380032 14492 380038 14544
rect 45186 14424 45192 14476
rect 45244 14464 45250 14476
rect 415394 14464 415400 14476
rect 45244 14436 415400 14464
rect 45244 14424 45250 14436
rect 415394 14424 415400 14436
rect 415452 14424 415458 14476
rect 166902 13336 166908 13388
rect 166960 13376 166966 13388
rect 295978 13376 295984 13388
rect 166960 13348 295984 13376
rect 166960 13336 166966 13348
rect 295978 13336 295984 13348
rect 296036 13336 296042 13388
rect 219250 13268 219256 13320
rect 219308 13308 219314 13320
rect 452838 13308 452844 13320
rect 219308 13280 452844 13308
rect 219308 13268 219314 13280
rect 452838 13268 452844 13280
rect 452896 13268 452902 13320
rect 83458 13200 83464 13252
rect 83516 13240 83522 13252
rect 355226 13240 355232 13252
rect 83516 13212 355232 13240
rect 83516 13200 83522 13212
rect 355226 13200 355232 13212
rect 355284 13200 355290 13252
rect 47670 13132 47676 13184
rect 47728 13172 47734 13184
rect 367002 13172 367008 13184
rect 47728 13144 367008 13172
rect 47728 13132 47734 13144
rect 367002 13132 367008 13144
rect 367060 13132 367066 13184
rect 381538 13132 381544 13184
rect 381596 13172 381602 13184
rect 446122 13172 446128 13184
rect 381596 13144 446128 13172
rect 381596 13132 381602 13144
rect 446122 13132 446128 13144
rect 446180 13132 446186 13184
rect 47854 13064 47860 13116
rect 47912 13104 47918 13116
rect 494698 13104 494704 13116
rect 47912 13076 494704 13104
rect 47912 13064 47918 13076
rect 494698 13064 494704 13076
rect 494756 13064 494762 13116
rect 208210 11976 208216 12028
rect 208268 12016 208274 12028
rect 446214 12016 446220 12028
rect 208268 11988 446220 12016
rect 208268 11976 208274 11988
rect 446214 11976 446220 11988
rect 446272 11976 446278 12028
rect 46566 11908 46572 11960
rect 46624 11948 46630 11960
rect 186130 11948 186136 11960
rect 46624 11920 186136 11948
rect 46624 11908 46630 11920
rect 186130 11908 186136 11920
rect 186188 11908 186194 11960
rect 190362 11908 190368 11960
rect 190420 11948 190426 11960
rect 452746 11948 452752 11960
rect 190420 11920 452752 11948
rect 190420 11908 190426 11920
rect 452746 11908 452752 11920
rect 452804 11908 452810 11960
rect 183462 11840 183468 11892
rect 183520 11880 183526 11892
rect 450354 11880 450360 11892
rect 183520 11852 450360 11880
rect 183520 11840 183526 11852
rect 450354 11840 450360 11852
rect 450412 11840 450418 11892
rect 126790 11772 126796 11824
rect 126848 11812 126854 11824
rect 450262 11812 450268 11824
rect 126848 11784 450268 11812
rect 126848 11772 126854 11784
rect 450262 11772 450268 11784
rect 450320 11772 450326 11824
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 445754 11744 445760 11756
rect 1360 11716 445760 11744
rect 1360 11704 1366 11716
rect 445754 11704 445760 11716
rect 445812 11704 445818 11756
rect 399846 11636 399852 11688
rect 399904 11676 399910 11688
rect 400122 11676 400128 11688
rect 399904 11648 400128 11676
rect 399904 11636 399910 11648
rect 400122 11636 400128 11648
rect 400180 11636 400186 11688
rect 423766 11636 423772 11688
rect 423824 11676 423830 11688
rect 424962 11676 424968 11688
rect 423824 11648 424968 11676
rect 423824 11636 423830 11648
rect 424962 11636 424968 11648
rect 425020 11636 425026 11688
rect 51902 10752 51908 10804
rect 51960 10792 51966 10804
rect 319714 10792 319720 10804
rect 51960 10764 319720 10792
rect 51960 10752 51966 10764
rect 319714 10752 319720 10764
rect 319772 10752 319778 10804
rect 125502 10684 125508 10736
rect 125560 10724 125566 10736
rect 448698 10724 448704 10736
rect 125560 10696 448704 10724
rect 125560 10684 125566 10696
rect 448698 10684 448704 10696
rect 448756 10684 448762 10736
rect 50614 10616 50620 10668
rect 50672 10656 50678 10668
rect 401318 10656 401324 10668
rect 50672 10628 401324 10656
rect 50672 10616 50678 10628
rect 401318 10616 401324 10628
rect 401376 10616 401382 10668
rect 50522 10548 50528 10600
rect 50580 10588 50586 10600
rect 411898 10588 411904 10600
rect 50580 10560 411904 10588
rect 50580 10548 50586 10560
rect 411898 10548 411904 10560
rect 411956 10548 411962 10600
rect 50430 10480 50436 10532
rect 50488 10520 50494 10532
rect 431954 10520 431960 10532
rect 50488 10492 431960 10520
rect 50488 10480 50494 10492
rect 431954 10480 431960 10492
rect 432012 10480 432018 10532
rect 50338 10412 50344 10464
rect 50396 10452 50402 10464
rect 449894 10452 449900 10464
rect 50396 10424 449900 10452
rect 50396 10412 50402 10424
rect 449894 10412 449900 10424
rect 449952 10412 449958 10464
rect 50890 10344 50896 10396
rect 50948 10384 50954 10396
rect 468386 10384 468392 10396
rect 50948 10356 468392 10384
rect 50948 10344 50954 10356
rect 468386 10344 468392 10356
rect 468444 10344 468450 10396
rect 50798 10276 50804 10328
rect 50856 10316 50862 10328
rect 479334 10316 479340 10328
rect 50856 10288 479340 10316
rect 50856 10276 50862 10288
rect 479334 10276 479340 10288
rect 479392 10276 479398 10328
rect 515398 10276 515404 10328
rect 515456 10316 515462 10328
rect 562042 10316 562048 10328
rect 515456 10288 562048 10316
rect 515456 10276 515462 10288
rect 562042 10276 562048 10288
rect 562100 10276 562106 10328
rect 222746 9596 222752 9648
rect 222804 9636 222810 9648
rect 440878 9636 440884 9648
rect 222804 9608 440884 9636
rect 222804 9596 222810 9608
rect 440878 9596 440884 9608
rect 440936 9596 440942 9648
rect 52362 9528 52368 9580
rect 52420 9568 52426 9580
rect 277118 9568 277124 9580
rect 52420 9540 277124 9568
rect 52420 9528 52426 9540
rect 277118 9528 277124 9540
rect 277176 9528 277182 9580
rect 52178 9460 52184 9512
rect 52236 9500 52242 9512
rect 280706 9500 280712 9512
rect 52236 9472 280712 9500
rect 52236 9460 52242 9472
rect 280706 9460 280712 9472
rect 280764 9460 280770 9512
rect 197906 9392 197912 9444
rect 197964 9432 197970 9444
rect 440326 9432 440332 9444
rect 197964 9404 440332 9432
rect 197964 9392 197970 9404
rect 440326 9392 440332 9404
rect 440384 9392 440390 9444
rect 53006 9324 53012 9376
rect 53064 9364 53070 9376
rect 304350 9364 304356 9376
rect 53064 9336 304356 9364
rect 53064 9324 53070 9336
rect 304350 9324 304356 9336
rect 304408 9324 304414 9376
rect 53466 9256 53472 9308
rect 53524 9296 53530 9308
rect 311434 9296 311440 9308
rect 53524 9268 311440 9296
rect 53524 9256 53530 9268
rect 311434 9256 311440 9268
rect 311492 9256 311498 9308
rect 51442 9188 51448 9240
rect 51500 9228 51506 9240
rect 312630 9228 312636 9240
rect 51500 9200 312636 9228
rect 51500 9188 51506 9200
rect 312630 9188 312636 9200
rect 312688 9188 312694 9240
rect 53190 9120 53196 9172
rect 53248 9160 53254 9172
rect 318518 9160 318524 9172
rect 53248 9132 318524 9160
rect 53248 9120 53254 9132
rect 318518 9120 318524 9132
rect 318576 9120 318582 9172
rect 320818 9120 320824 9172
rect 320876 9160 320882 9172
rect 348050 9160 348056 9172
rect 320876 9132 348056 9160
rect 320876 9120 320882 9132
rect 348050 9120 348056 9132
rect 348108 9120 348114 9172
rect 53558 9052 53564 9104
rect 53616 9092 53622 9104
rect 346946 9092 346952 9104
rect 53616 9064 346952 9092
rect 53616 9052 53622 9064
rect 346946 9052 346952 9064
rect 347004 9052 347010 9104
rect 53742 8984 53748 9036
rect 53800 9024 53806 9036
rect 378870 9024 378876 9036
rect 53800 8996 378876 9024
rect 53800 8984 53806 8996
rect 378870 8984 378876 8996
rect 378928 8984 378934 9036
rect 51718 8916 51724 8968
rect 51776 8956 51782 8968
rect 571518 8956 571524 8968
rect 51776 8928 571524 8956
rect 51776 8916 51782 8928
rect 571518 8916 571524 8928
rect 571576 8916 571582 8968
rect 52270 8848 52276 8900
rect 52328 8888 52334 8900
rect 270034 8888 270040 8900
rect 52328 8860 270040 8888
rect 52328 8848 52334 8860
rect 270034 8848 270040 8860
rect 270092 8848 270098 8900
rect 51626 8780 51632 8832
rect 51684 8820 51690 8832
rect 266538 8820 266544 8832
rect 51684 8792 266544 8820
rect 51684 8780 51690 8792
rect 266538 8780 266544 8792
rect 266596 8780 266602 8832
rect 53282 8712 53288 8764
rect 53340 8752 53346 8764
rect 268838 8752 268844 8764
rect 53340 8724 268844 8752
rect 53340 8712 53346 8724
rect 268838 8712 268844 8724
rect 268896 8712 268902 8764
rect 252370 8644 252376 8696
rect 252428 8684 252434 8696
rect 447870 8684 447876 8696
rect 252428 8656 447876 8684
rect 252428 8644 252434 8656
rect 447870 8644 447876 8656
rect 447928 8644 447934 8696
rect 262950 8576 262956 8628
rect 263008 8616 263014 8628
rect 447410 8616 447416 8628
rect 263008 8588 447416 8616
rect 263008 8576 263014 8588
rect 447410 8576 447416 8588
rect 447468 8576 447474 8628
rect 265342 8508 265348 8560
rect 265400 8548 265406 8560
rect 443638 8548 443644 8560
rect 265400 8520 443644 8548
rect 265400 8508 265406 8520
rect 443638 8508 443644 8520
rect 443696 8508 443702 8560
rect 259454 8440 259460 8492
rect 259512 8480 259518 8492
rect 383654 8480 383660 8492
rect 259512 8452 383660 8480
rect 259512 8440 259518 8452
rect 383654 8440 383660 8452
rect 383712 8440 383718 8492
rect 50982 8236 50988 8288
rect 51040 8276 51046 8288
rect 160186 8276 160192 8288
rect 51040 8248 160192 8276
rect 51040 8236 51046 8248
rect 160186 8236 160192 8248
rect 160244 8236 160250 8288
rect 169570 8236 169576 8288
rect 169628 8276 169634 8288
rect 440418 8276 440424 8288
rect 169628 8248 440424 8276
rect 169628 8236 169634 8248
rect 440418 8236 440424 8248
rect 440476 8236 440482 8288
rect 147122 8168 147128 8220
rect 147180 8208 147186 8220
rect 443454 8208 443460 8220
rect 147180 8180 443460 8208
rect 147180 8168 147186 8180
rect 443454 8168 443460 8180
rect 443512 8168 443518 8220
rect 54570 8100 54576 8152
rect 54628 8140 54634 8152
rect 194410 8140 194416 8152
rect 54628 8112 194416 8140
rect 54628 8100 54634 8112
rect 194410 8100 194416 8112
rect 194468 8100 194474 8152
rect 219342 8100 219348 8152
rect 219400 8140 219406 8152
rect 545482 8140 545488 8152
rect 219400 8112 545488 8140
rect 219400 8100 219406 8112
rect 545482 8100 545488 8112
rect 545540 8100 545546 8152
rect 55858 8032 55864 8084
rect 55916 8072 55922 8084
rect 434438 8072 434444 8084
rect 55916 8044 434444 8072
rect 55916 8032 55922 8044
rect 434438 8032 434444 8044
rect 434496 8032 434502 8084
rect 56134 7964 56140 8016
rect 56192 8004 56198 8016
rect 437934 8004 437940 8016
rect 56192 7976 437940 8004
rect 56192 7964 56198 7976
rect 437934 7964 437940 7976
rect 437992 7964 437998 8016
rect 126882 7896 126888 7948
rect 126940 7936 126946 7948
rect 517146 7936 517152 7948
rect 126940 7908 517152 7936
rect 126940 7896 126946 7908
rect 517146 7896 517152 7908
rect 517204 7896 517210 7948
rect 55766 7828 55772 7880
rect 55824 7868 55830 7880
rect 466270 7868 466276 7880
rect 55824 7840 466276 7868
rect 55824 7828 55830 7840
rect 466270 7828 466276 7840
rect 466328 7828 466334 7880
rect 56410 7760 56416 7812
rect 56468 7800 56474 7812
rect 469858 7800 469864 7812
rect 56468 7772 469864 7800
rect 56468 7760 56474 7772
rect 469858 7760 469864 7772
rect 469916 7760 469922 7812
rect 54110 7692 54116 7744
rect 54168 7732 54174 7744
rect 549070 7732 549076 7744
rect 54168 7704 549076 7732
rect 54168 7692 54174 7704
rect 549070 7692 549076 7704
rect 549128 7692 549134 7744
rect 53926 7624 53932 7676
rect 53984 7664 53990 7676
rect 566826 7664 566832 7676
rect 53984 7636 566832 7664
rect 53984 7624 53990 7636
rect 566826 7624 566832 7636
rect 566884 7624 566890 7676
rect 54386 7556 54392 7608
rect 54444 7596 54450 7608
rect 577406 7596 577412 7608
rect 54444 7568 577412 7596
rect 54444 7556 54450 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 173158 7488 173164 7540
rect 173216 7528 173222 7540
rect 440970 7528 440976 7540
rect 173216 7500 440976 7528
rect 173216 7488 173222 7500
rect 440970 7488 440976 7500
rect 441028 7488 441034 7540
rect 227530 7420 227536 7472
rect 227588 7460 227594 7472
rect 459186 7460 459192 7472
rect 227588 7432 459192 7460
rect 227588 7420 227594 7432
rect 459186 7420 459192 7432
rect 459244 7420 459250 7472
rect 147582 7352 147588 7404
rect 147640 7392 147646 7404
rect 342070 7392 342076 7404
rect 147640 7364 342076 7392
rect 147640 7352 147646 7364
rect 342070 7352 342076 7364
rect 342128 7352 342134 7404
rect 51350 7284 51356 7336
rect 51408 7324 51414 7336
rect 234706 7324 234712 7336
rect 51408 7296 234712 7324
rect 51408 7284 51414 7296
rect 234706 7284 234712 7296
rect 234764 7284 234770 7336
rect 263502 7284 263508 7336
rect 263560 7324 263566 7336
rect 395338 7324 395344 7336
rect 263560 7296 395344 7324
rect 263560 7284 263566 7296
rect 395338 7284 395344 7296
rect 395396 7284 395402 7336
rect 224770 7216 224776 7268
rect 224828 7256 224834 7268
rect 391842 7256 391848 7268
rect 224828 7228 391848 7256
rect 224828 7216 224834 7228
rect 391842 7216 391848 7228
rect 391900 7216 391906 7268
rect 203886 7148 203892 7200
rect 203944 7188 203950 7200
rect 336826 7188 336832 7200
rect 203944 7160 336832 7188
rect 203944 7148 203950 7160
rect 336826 7148 336832 7160
rect 336884 7148 336890 7200
rect 228726 7080 228732 7132
rect 228784 7120 228790 7132
rect 358906 7120 358912 7132
rect 228784 7092 358912 7120
rect 228784 7080 228790 7092
rect 358906 7080 358912 7092
rect 358964 7080 358970 7132
rect 199930 7012 199936 7064
rect 199988 7052 199994 7064
rect 241698 7052 241704 7064
rect 199988 7024 241704 7052
rect 199988 7012 199994 7024
rect 241698 7012 241704 7024
rect 241756 7012 241762 7064
rect 266262 7012 266268 7064
rect 266320 7052 266326 7064
rect 388254 7052 388260 7064
rect 266320 7024 388260 7052
rect 266320 7012 266326 7024
rect 388254 7012 388260 7024
rect 388312 7012 388318 7064
rect 257890 6944 257896 6996
rect 257948 6984 257954 6996
rect 320910 6984 320916 6996
rect 257948 6956 320916 6984
rect 257948 6944 257954 6956
rect 320910 6944 320916 6956
rect 320968 6944 320974 6996
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 39298 6848 39304 6860
rect 3476 6820 39304 6848
rect 3476 6808 3482 6820
rect 39298 6808 39304 6820
rect 39356 6808 39362 6860
rect 69106 6808 69112 6860
rect 69164 6848 69170 6860
rect 350534 6848 350540 6860
rect 69164 6820 350540 6848
rect 69164 6808 69170 6820
rect 350534 6808 350540 6820
rect 350592 6808 350598 6860
rect 461670 6808 461676 6860
rect 461728 6848 461734 6860
rect 580166 6848 580172 6860
rect 461728 6820 580172 6848
rect 461728 6808 461734 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 54294 6740 54300 6792
rect 54352 6780 54358 6792
rect 176746 6780 176752 6792
rect 54352 6752 176752 6780
rect 54352 6740 54358 6752
rect 176746 6740 176752 6752
rect 176804 6740 176810 6792
rect 177942 6740 177948 6792
rect 178000 6780 178006 6792
rect 461578 6780 461584 6792
rect 178000 6752 461584 6780
rect 178000 6740 178006 6752
rect 461578 6740 461584 6752
rect 461636 6740 461642 6792
rect 116394 6672 116400 6724
rect 116452 6712 116458 6724
rect 448882 6712 448888 6724
rect 116452 6684 448888 6712
rect 116452 6672 116458 6684
rect 448882 6672 448888 6684
rect 448940 6672 448946 6724
rect 90358 6604 90364 6656
rect 90416 6644 90422 6656
rect 427814 6644 427820 6656
rect 90416 6616 427820 6644
rect 90416 6604 90422 6616
rect 427814 6604 427820 6616
rect 427872 6604 427878 6656
rect 55122 6536 55128 6588
rect 55180 6576 55186 6588
rect 187326 6576 187332 6588
rect 55180 6548 187332 6576
rect 55180 6536 55186 6548
rect 187326 6536 187332 6548
rect 187384 6536 187390 6588
rect 195882 6536 195888 6588
rect 195940 6576 195946 6588
rect 580994 6576 581000 6588
rect 195940 6548 581000 6576
rect 195940 6536 195946 6548
rect 580994 6536 581000 6548
rect 581052 6536 581058 6588
rect 18230 6468 18236 6520
rect 18288 6508 18294 6520
rect 416866 6508 416872 6520
rect 18288 6480 416872 6508
rect 18288 6468 18294 6480
rect 416866 6468 416872 6480
rect 416924 6468 416930 6520
rect 427262 6468 427268 6520
rect 427320 6508 427326 6520
rect 454126 6508 454132 6520
rect 427320 6480 454132 6508
rect 427320 6468 427326 6480
rect 454126 6468 454132 6480
rect 454184 6468 454190 6520
rect 50154 6400 50160 6452
rect 50212 6440 50218 6452
rect 448974 6440 448980 6452
rect 50212 6412 448980 6440
rect 50212 6400 50218 6412
rect 448974 6400 448980 6412
rect 449032 6400 449038 6452
rect 41874 6332 41880 6384
rect 41932 6372 41938 6384
rect 448514 6372 448520 6384
rect 41932 6344 448520 6372
rect 41932 6332 41938 6344
rect 448514 6332 448520 6344
rect 448572 6332 448578 6384
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 449158 6304 449164 6316
rect 19484 6276 449164 6304
rect 19484 6264 19490 6276
rect 449158 6264 449164 6276
rect 449216 6264 449222 6316
rect 54938 6196 54944 6248
rect 54996 6236 55002 6248
rect 69658 6236 69664 6248
rect 54996 6208 69664 6236
rect 54996 6196 55002 6208
rect 69658 6196 69664 6208
rect 69716 6196 69722 6248
rect 74442 6196 74448 6248
rect 74500 6236 74506 6248
rect 515950 6236 515956 6248
rect 74500 6208 515956 6236
rect 74500 6196 74506 6208
rect 515950 6196 515956 6208
rect 516008 6196 516014 6248
rect 58894 6128 58900 6180
rect 58952 6168 58958 6180
rect 523034 6168 523040 6180
rect 58952 6140 523040 6168
rect 58952 6128 58958 6140
rect 523034 6128 523040 6140
rect 523092 6128 523098 6180
rect 31294 6060 31300 6112
rect 31352 6100 31358 6112
rect 273254 6100 273260 6112
rect 31352 6072 273260 6100
rect 31352 6060 31358 6072
rect 273254 6060 273260 6072
rect 273312 6060 273318 6112
rect 301958 6060 301964 6112
rect 302016 6100 302022 6112
rect 447226 6100 447232 6112
rect 302016 6072 447232 6100
rect 302016 6060 302022 6072
rect 447226 6060 447232 6072
rect 447284 6060 447290 6112
rect 86862 5992 86868 6044
rect 86920 6032 86926 6044
rect 317414 6032 317420 6044
rect 86920 6004 317420 6032
rect 86920 5992 86926 6004
rect 317414 5992 317420 6004
rect 317472 5992 317478 6044
rect 322106 5992 322112 6044
rect 322164 6032 322170 6044
rect 444466 6032 444472 6044
rect 322164 6004 444472 6032
rect 322164 5992 322170 6004
rect 444466 5992 444472 6004
rect 444524 5992 444530 6044
rect 101030 5924 101036 5976
rect 101088 5964 101094 5976
rect 306374 5964 306380 5976
rect 101088 5936 306380 5964
rect 101088 5924 101094 5936
rect 306374 5924 306380 5936
rect 306432 5924 306438 5976
rect 330386 5924 330392 5976
rect 330444 5964 330450 5976
rect 447318 5964 447324 5976
rect 330444 5936 447324 5964
rect 330444 5924 330450 5936
rect 447318 5924 447324 5936
rect 447376 5924 447382 5976
rect 114002 5856 114008 5908
rect 114060 5896 114066 5908
rect 289814 5896 289820 5908
rect 114060 5868 289820 5896
rect 114060 5856 114066 5868
rect 289814 5856 289820 5868
rect 289872 5856 289878 5908
rect 59538 5788 59544 5840
rect 59596 5828 59602 5840
rect 153010 5828 153016 5840
rect 59596 5800 153016 5828
rect 59596 5788 59602 5800
rect 153010 5788 153016 5800
rect 153068 5788 153074 5840
rect 112990 5448 112996 5500
rect 113048 5488 113054 5500
rect 317322 5488 317328 5500
rect 113048 5460 317328 5488
rect 113048 5448 113054 5460
rect 317322 5448 317328 5460
rect 317380 5448 317386 5500
rect 356330 5448 356336 5500
rect 356388 5488 356394 5500
rect 422386 5488 422392 5500
rect 356388 5460 422392 5488
rect 356388 5448 356394 5460
rect 422386 5448 422392 5460
rect 422444 5448 422450 5500
rect 53650 5380 53656 5432
rect 53708 5420 53714 5432
rect 151814 5420 151820 5432
rect 53708 5392 151820 5420
rect 53708 5380 53714 5392
rect 151814 5380 151820 5392
rect 151872 5380 151878 5432
rect 225138 5380 225144 5432
rect 225196 5420 225202 5432
rect 443086 5420 443092 5432
rect 225196 5392 443092 5420
rect 225196 5380 225202 5392
rect 443086 5380 443092 5392
rect 443144 5380 443150 5432
rect 59354 5312 59360 5364
rect 59412 5352 59418 5364
rect 306742 5352 306748 5364
rect 59412 5324 306748 5352
rect 59412 5312 59418 5324
rect 306742 5312 306748 5324
rect 306800 5312 306806 5364
rect 316218 5312 316224 5364
rect 316276 5352 316282 5364
rect 447134 5352 447140 5364
rect 316276 5324 447140 5352
rect 316276 5312 316282 5324
rect 447134 5312 447140 5324
rect 447192 5312 447198 5364
rect 59170 5244 59176 5296
rect 59228 5284 59234 5296
rect 196802 5284 196808 5296
rect 59228 5256 196808 5284
rect 59228 5244 59234 5256
rect 196802 5244 196808 5256
rect 196860 5244 196866 5296
rect 208302 5244 208308 5296
rect 208360 5284 208366 5296
rect 455690 5284 455696 5296
rect 208360 5256 455696 5284
rect 208360 5244 208366 5256
rect 455690 5244 455696 5256
rect 455748 5244 455754 5296
rect 58802 5176 58808 5228
rect 58860 5216 58866 5228
rect 164878 5216 164884 5228
rect 58860 5188 164884 5216
rect 58860 5176 58866 5188
rect 164878 5176 164884 5188
rect 164936 5176 164942 5228
rect 171962 5176 171968 5228
rect 172020 5216 172026 5228
rect 430574 5216 430580 5228
rect 172020 5188 430580 5216
rect 172020 5176 172026 5188
rect 430574 5176 430580 5188
rect 430632 5176 430638 5228
rect 132954 5108 132960 5160
rect 133012 5148 133018 5160
rect 391934 5148 391940 5160
rect 133012 5120 391940 5148
rect 133012 5108 133018 5120
rect 391934 5108 391940 5120
rect 391992 5108 391998 5160
rect 394234 5108 394240 5160
rect 394292 5148 394298 5160
rect 440142 5148 440148 5160
rect 394292 5120 440148 5148
rect 394292 5108 394298 5120
rect 440142 5108 440148 5120
rect 440200 5108 440206 5160
rect 63310 5040 63316 5092
rect 63368 5080 63374 5092
rect 324406 5080 324412 5092
rect 63368 5052 324412 5080
rect 63368 5040 63374 5052
rect 324406 5040 324412 5052
rect 324464 5040 324470 5092
rect 335078 5040 335084 5092
rect 335136 5080 335142 5092
rect 425054 5080 425060 5092
rect 335136 5052 425060 5080
rect 335136 5040 335142 5052
rect 425054 5040 425060 5052
rect 425112 5040 425118 5092
rect 426158 5040 426164 5092
rect 426216 5080 426222 5092
rect 447686 5080 447692 5092
rect 426216 5052 447692 5080
rect 426216 5040 426222 5052
rect 447686 5040 447692 5052
rect 447744 5040 447750 5092
rect 66070 4972 66076 5024
rect 66128 5012 66134 5024
rect 358630 5012 358636 5024
rect 66128 4984 358636 5012
rect 66128 4972 66134 4984
rect 358630 4972 358636 4984
rect 358688 4972 358694 5024
rect 388441 5015 388499 5021
rect 388441 4981 388453 5015
rect 388487 5012 388499 5015
rect 572714 5012 572720 5024
rect 388487 4984 572720 5012
rect 388487 4981 388499 4984
rect 388441 4975 388499 4981
rect 572714 4972 572720 4984
rect 572772 4972 572778 5024
rect 17034 4904 17040 4956
rect 17092 4944 17098 4956
rect 234614 4944 234620 4956
rect 17092 4916 234620 4944
rect 17092 4904 17098 4916
rect 234614 4904 234620 4916
rect 234672 4904 234678 4956
rect 244182 4904 244188 4956
rect 244240 4944 244246 4956
rect 537202 4944 537208 4956
rect 244240 4916 537208 4944
rect 244240 4904 244246 4916
rect 537202 4904 537208 4916
rect 537260 4904 537266 4956
rect 50706 4836 50712 4888
rect 50764 4876 50770 4888
rect 156598 4876 156604 4888
rect 50764 4848 156604 4876
rect 50764 4836 50770 4848
rect 156598 4836 156604 4848
rect 156656 4836 156662 4888
rect 161382 4836 161388 4888
rect 161440 4876 161446 4888
rect 533706 4876 533712 4888
rect 161440 4848 533712 4876
rect 161440 4836 161446 4848
rect 533706 4836 533712 4848
rect 533764 4836 533770 4888
rect 537478 4836 537484 4888
rect 537536 4876 537542 4888
rect 538398 4876 538404 4888
rect 537536 4848 538404 4876
rect 537536 4836 537542 4848
rect 538398 4836 538404 4848
rect 538456 4836 538462 4888
rect 56502 4768 56508 4820
rect 56560 4808 56566 4820
rect 448514 4808 448520 4820
rect 56560 4780 448520 4808
rect 56560 4768 56566 4780
rect 448514 4768 448520 4780
rect 448572 4768 448578 4820
rect 511258 4768 511264 4820
rect 511316 4808 511322 4820
rect 520734 4808 520740 4820
rect 511316 4780 520740 4808
rect 511316 4768 511322 4780
rect 520734 4768 520740 4780
rect 520792 4768 520798 4820
rect 68922 4700 68928 4752
rect 68980 4740 68986 4752
rect 264146 4740 264152 4752
rect 68980 4712 264152 4740
rect 68980 4700 68986 4712
rect 264146 4700 264152 4712
rect 264204 4700 264210 4752
rect 274818 4700 274824 4752
rect 274876 4740 274882 4752
rect 274876 4712 441614 4740
rect 274876 4700 274882 4712
rect 59446 4632 59452 4684
rect 59504 4672 59510 4684
rect 249978 4672 249984 4684
rect 59504 4644 249984 4672
rect 59504 4632 59510 4644
rect 249978 4632 249984 4644
rect 250036 4632 250042 4684
rect 260650 4632 260656 4684
rect 260708 4672 260714 4684
rect 441586 4672 441614 4712
rect 443270 4672 443276 4684
rect 260708 4644 436784 4672
rect 441586 4644 443276 4672
rect 260708 4632 260714 4644
rect 51810 4564 51816 4616
rect 51868 4604 51874 4616
rect 142430 4604 142436 4616
rect 51868 4576 142436 4604
rect 51868 4564 51874 4576
rect 142430 4564 142436 4576
rect 142488 4564 142494 4616
rect 146202 4564 146208 4616
rect 146260 4604 146266 4616
rect 267734 4604 267740 4616
rect 146260 4576 267740 4604
rect 146260 4564 146266 4576
rect 267734 4564 267740 4576
rect 267792 4564 267798 4616
rect 278314 4564 278320 4616
rect 278372 4604 278378 4616
rect 436756 4604 436784 4644
rect 443270 4632 443276 4644
rect 443328 4632 443334 4684
rect 278372 4576 435772 4604
rect 436756 4576 441614 4604
rect 278372 4564 278378 4576
rect 52914 4496 52920 4548
rect 52972 4536 52978 4548
rect 141234 4536 141240 4548
rect 52972 4508 141240 4536
rect 52972 4496 52978 4508
rect 141234 4496 141240 4508
rect 141292 4496 141298 4548
rect 143442 4496 143448 4548
rect 143500 4536 143506 4548
rect 299658 4536 299664 4548
rect 143500 4508 299664 4536
rect 143500 4496 143506 4508
rect 299658 4496 299664 4508
rect 299716 4496 299722 4548
rect 313826 4496 313832 4548
rect 313884 4536 313890 4548
rect 435744 4536 435772 4576
rect 439498 4536 439504 4548
rect 313884 4508 432092 4536
rect 435744 4508 439504 4536
rect 313884 4496 313890 4508
rect 58710 4428 58716 4480
rect 58768 4468 58774 4480
rect 136450 4468 136456 4480
rect 58768 4440 136456 4468
rect 58768 4428 58774 4440
rect 136450 4428 136456 4440
rect 136508 4428 136514 4480
rect 140038 4428 140044 4480
rect 140096 4468 140102 4480
rect 204254 4468 204260 4480
rect 140096 4440 204260 4468
rect 140096 4428 140102 4440
rect 204254 4428 204260 4440
rect 204312 4428 204318 4480
rect 239306 4428 239312 4480
rect 239364 4468 239370 4480
rect 364426 4468 364432 4480
rect 239364 4440 364432 4468
rect 239364 4428 239370 4440
rect 364426 4428 364432 4440
rect 364484 4428 364490 4480
rect 379422 4428 379428 4480
rect 379480 4468 379486 4480
rect 388441 4471 388499 4477
rect 388441 4468 388453 4471
rect 379480 4440 388453 4468
rect 379480 4428 379486 4440
rect 388441 4437 388453 4440
rect 388487 4437 388499 4471
rect 388441 4431 388499 4437
rect 413094 4428 413100 4480
rect 413152 4468 413158 4480
rect 413152 4440 431954 4468
rect 413152 4428 413158 4440
rect 169662 4360 169668 4412
rect 169720 4400 169726 4412
rect 271230 4400 271236 4412
rect 169720 4372 271236 4400
rect 169720 4360 169726 4372
rect 271230 4360 271236 4372
rect 271288 4360 271294 4412
rect 298738 4360 298744 4412
rect 298796 4400 298802 4412
rect 397730 4400 397736 4412
rect 298796 4372 397736 4400
rect 298796 4360 298802 4372
rect 397730 4360 397736 4372
rect 397788 4360 397794 4412
rect 234430 4292 234436 4344
rect 234488 4332 234494 4344
rect 242894 4332 242900 4344
rect 234488 4304 242900 4332
rect 234488 4292 234494 4304
rect 242894 4292 242900 4304
rect 242952 4292 242958 4344
rect 292574 4292 292580 4344
rect 292632 4332 292638 4344
rect 339494 4332 339500 4344
rect 292632 4304 339500 4332
rect 292632 4292 292638 4304
rect 339494 4292 339500 4304
rect 339552 4292 339558 4344
rect 431926 4332 431954 4440
rect 432064 4400 432092 4508
rect 439498 4496 439504 4508
rect 439556 4496 439562 4548
rect 441586 4536 441614 4576
rect 443362 4536 443368 4548
rect 441586 4508 443368 4536
rect 443362 4496 443368 4508
rect 443420 4496 443426 4548
rect 460198 4496 460204 4548
rect 460256 4536 460262 4548
rect 462774 4536 462780 4548
rect 460256 4508 462780 4536
rect 460256 4496 460262 4508
rect 462774 4496 462780 4508
rect 462832 4496 462838 4548
rect 475378 4496 475384 4548
rect 475436 4536 475442 4548
rect 481726 4536 481732 4548
rect 475436 4508 481732 4536
rect 475436 4496 475442 4508
rect 481726 4496 481732 4508
rect 481784 4496 481790 4548
rect 443730 4400 443736 4412
rect 432064 4372 443736 4400
rect 443730 4360 443736 4372
rect 443788 4360 443794 4412
rect 440602 4332 440608 4344
rect 431926 4304 440608 4332
rect 440602 4292 440608 4304
rect 440660 4292 440666 4344
rect 327994 4224 328000 4276
rect 328052 4264 328058 4276
rect 372706 4264 372712 4276
rect 328052 4236 372712 4264
rect 328052 4224 328058 4236
rect 372706 4224 372712 4236
rect 372764 4224 372770 4276
rect 160094 4156 160100 4208
rect 160152 4196 160158 4208
rect 161290 4196 161296 4208
rect 160152 4168 161296 4196
rect 160152 4156 160158 4168
rect 161290 4156 161296 4168
rect 161348 4156 161354 4208
rect 407758 4156 407764 4208
rect 407816 4196 407822 4208
rect 409598 4196 409604 4208
rect 407816 4168 409604 4196
rect 407816 4156 407822 4168
rect 409598 4156 409604 4168
rect 409656 4156 409662 4208
rect 445018 4156 445024 4208
rect 445076 4196 445082 4208
rect 449986 4196 449992 4208
rect 445076 4168 449992 4196
rect 445076 4156 445082 4168
rect 449986 4156 449992 4168
rect 450044 4156 450050 4208
rect 533338 4156 533344 4208
rect 533396 4196 533402 4208
rect 534902 4196 534908 4208
rect 533396 4168 534908 4196
rect 533396 4156 533402 4168
rect 534902 4156 534908 4168
rect 534960 4156 534966 4208
rect 57054 4088 57060 4140
rect 57112 4128 57118 4140
rect 71498 4128 71504 4140
rect 57112 4100 71504 4128
rect 57112 4088 57118 4100
rect 71498 4088 71504 4100
rect 71556 4088 71562 4140
rect 71682 4088 71688 4140
rect 71740 4128 71746 4140
rect 71740 4100 72740 4128
rect 71740 4088 71746 4100
rect 57882 4020 57888 4072
rect 57940 4060 57946 4072
rect 72602 4060 72608 4072
rect 57940 4032 72608 4060
rect 57940 4020 57946 4032
rect 72602 4020 72608 4032
rect 72660 4020 72666 4072
rect 72712 4060 72740 4100
rect 76190 4088 76196 4140
rect 76248 4128 76254 4140
rect 77202 4128 77208 4140
rect 76248 4100 77208 4128
rect 76248 4088 76254 4100
rect 77202 4088 77208 4100
rect 77260 4088 77266 4140
rect 77297 4131 77355 4137
rect 77297 4097 77309 4131
rect 77343 4128 77355 4131
rect 442166 4128 442172 4140
rect 77343 4100 442172 4128
rect 77343 4097 77355 4100
rect 77297 4091 77355 4097
rect 442166 4088 442172 4100
rect 442224 4088 442230 4140
rect 536098 4088 536104 4140
rect 536156 4128 536162 4140
rect 539594 4128 539600 4140
rect 536156 4100 539600 4128
rect 536156 4088 536162 4100
rect 539594 4088 539600 4100
rect 539652 4088 539658 4140
rect 441614 4060 441620 4072
rect 72712 4032 441620 4060
rect 441614 4020 441620 4032
rect 441672 4020 441678 4072
rect 485038 4020 485044 4072
rect 485096 4060 485102 4072
rect 492306 4060 492312 4072
rect 485096 4032 492312 4060
rect 485096 4020 485102 4032
rect 492306 4020 492312 4032
rect 492364 4020 492370 4072
rect 529198 4020 529204 4072
rect 529256 4060 529262 4072
rect 546678 4060 546684 4072
rect 529256 4032 546684 4060
rect 529256 4020 529262 4032
rect 546678 4020 546684 4032
rect 546736 4020 546742 4072
rect 64846 3964 66300 3992
rect 53742 3884 53748 3936
rect 53800 3924 53806 3936
rect 64846 3924 64874 3964
rect 53800 3896 64874 3924
rect 53800 3884 53806 3896
rect 65518 3884 65524 3936
rect 65576 3924 65582 3936
rect 66162 3924 66168 3936
rect 65576 3896 66168 3924
rect 65576 3884 65582 3896
rect 66162 3884 66168 3896
rect 66220 3884 66226 3936
rect 66272 3924 66300 3964
rect 70302 3952 70308 4004
rect 70360 3992 70366 4004
rect 311894 3992 311900 4004
rect 70360 3964 311900 3992
rect 70360 3952 70366 3964
rect 311894 3952 311900 3964
rect 311952 3952 311958 4004
rect 340966 3952 340972 4004
rect 341024 3992 341030 4004
rect 342162 3992 342168 4004
rect 341024 3964 342168 3992
rect 341024 3952 341030 3964
rect 342162 3952 342168 3964
rect 342220 3952 342226 4004
rect 440326 3952 440332 4004
rect 440384 3992 440390 4004
rect 455414 3992 455420 4004
rect 440384 3964 455420 3992
rect 440384 3952 440390 3964
rect 455414 3952 455420 3964
rect 455472 3952 455478 4004
rect 520918 3952 520924 4004
rect 520976 3992 520982 4004
rect 524325 3995 524383 4001
rect 524325 3992 524337 3995
rect 520976 3964 524337 3992
rect 520976 3952 520982 3964
rect 524325 3961 524337 3964
rect 524371 3961 524383 3995
rect 524325 3955 524383 3961
rect 531958 3952 531964 4004
rect 532016 3992 532022 4004
rect 553762 3992 553768 4004
rect 532016 3964 553768 3992
rect 532016 3952 532022 3964
rect 553762 3952 553768 3964
rect 553820 3952 553826 4004
rect 70394 3924 70400 3936
rect 66272 3896 70400 3924
rect 70394 3884 70400 3896
rect 70452 3884 70458 3936
rect 71590 3884 71596 3936
rect 71648 3924 71654 3936
rect 77297 3927 77355 3933
rect 77297 3924 77309 3927
rect 71648 3896 77309 3924
rect 71648 3884 71654 3896
rect 77297 3893 77309 3896
rect 77343 3893 77355 3927
rect 77297 3887 77355 3893
rect 78582 3884 78588 3936
rect 78640 3924 78646 3936
rect 347774 3924 347780 3936
rect 78640 3896 347780 3924
rect 78640 3884 78646 3896
rect 347774 3884 347780 3896
rect 347832 3884 347838 3936
rect 418982 3884 418988 3936
rect 419040 3924 419046 3936
rect 441890 3924 441896 3936
rect 419040 3896 441896 3924
rect 419040 3884 419046 3896
rect 441890 3884 441896 3896
rect 441948 3884 441954 3936
rect 523678 3884 523684 3936
rect 523736 3924 523742 3936
rect 536098 3924 536104 3936
rect 523736 3896 536104 3924
rect 523736 3884 523742 3896
rect 536098 3884 536104 3896
rect 536156 3884 536162 3936
rect 538858 3884 538864 3936
rect 538916 3924 538922 3936
rect 564434 3924 564440 3936
rect 538916 3896 564440 3924
rect 538916 3884 538922 3896
rect 564434 3884 564440 3896
rect 564492 3884 564498 3936
rect 39574 3816 39580 3868
rect 39632 3856 39638 3868
rect 307757 3859 307815 3865
rect 307757 3856 307769 3859
rect 39632 3828 307769 3856
rect 39632 3816 39638 3828
rect 307757 3825 307769 3828
rect 307803 3825 307815 3859
rect 307757 3819 307815 3825
rect 307846 3816 307852 3868
rect 307904 3856 307910 3868
rect 309042 3856 309048 3868
rect 307904 3828 309048 3856
rect 307904 3816 307910 3828
rect 309042 3816 309048 3828
rect 309100 3816 309106 3868
rect 324130 3816 324136 3868
rect 324188 3856 324194 3868
rect 454494 3856 454500 3868
rect 324188 3828 454500 3856
rect 324188 3816 324194 3828
rect 454494 3816 454500 3828
rect 454552 3816 454558 3868
rect 500218 3816 500224 3868
rect 500276 3856 500282 3868
rect 506474 3856 506480 3868
rect 500276 3828 506480 3856
rect 500276 3816 500282 3828
rect 506474 3816 506480 3828
rect 506532 3816 506538 3868
rect 518158 3816 518164 3868
rect 518216 3856 518222 3868
rect 532510 3856 532516 3868
rect 518216 3828 532516 3856
rect 518216 3816 518222 3828
rect 532510 3816 532516 3828
rect 532568 3816 532574 3868
rect 542998 3816 543004 3868
rect 543056 3856 543062 3868
rect 575106 3856 575112 3868
rect 543056 3828 575112 3856
rect 543056 3816 543062 3828
rect 575106 3816 575112 3828
rect 575164 3816 575170 3868
rect 56870 3748 56876 3800
rect 56928 3788 56934 3800
rect 102226 3788 102232 3800
rect 56928 3760 102232 3788
rect 56928 3748 56934 3760
rect 102226 3748 102232 3760
rect 102284 3748 102290 3800
rect 122282 3748 122288 3800
rect 122340 3788 122346 3800
rect 122742 3788 122748 3800
rect 122340 3760 122748 3788
rect 122340 3748 122346 3760
rect 122742 3748 122748 3760
rect 122800 3748 122806 3800
rect 127621 3791 127679 3797
rect 127621 3757 127633 3791
rect 127667 3788 127679 3791
rect 442350 3788 442356 3800
rect 127667 3760 442356 3788
rect 127667 3757 127679 3760
rect 127621 3751 127679 3757
rect 442350 3748 442356 3760
rect 442408 3748 442414 3800
rect 493318 3748 493324 3800
rect 493376 3788 493382 3800
rect 511258 3788 511264 3800
rect 493376 3760 511264 3788
rect 493376 3748 493382 3760
rect 511258 3748 511264 3760
rect 511316 3748 511322 3800
rect 518250 3748 518256 3800
rect 518308 3788 518314 3800
rect 521838 3788 521844 3800
rect 518308 3760 521844 3788
rect 518308 3748 518314 3760
rect 521838 3748 521844 3760
rect 521896 3748 521902 3800
rect 527910 3748 527916 3800
rect 527968 3788 527974 3800
rect 543182 3788 543188 3800
rect 527968 3760 543188 3788
rect 527968 3748 527974 3760
rect 543182 3748 543188 3760
rect 543240 3748 543246 3800
rect 545758 3748 545764 3800
rect 545816 3788 545822 3800
rect 578602 3788 578608 3800
rect 545816 3760 578608 3788
rect 545816 3748 545822 3760
rect 578602 3748 578608 3760
rect 578660 3748 578666 3800
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 361574 3720 361580 3732
rect 20680 3692 361580 3720
rect 20680 3680 20686 3692
rect 361574 3680 361580 3692
rect 361632 3680 361638 3732
rect 415486 3680 415492 3732
rect 415544 3720 415550 3732
rect 442626 3720 442632 3732
rect 415544 3692 442632 3720
rect 415544 3680 415550 3692
rect 442626 3680 442632 3692
rect 442684 3680 442690 3732
rect 494790 3680 494796 3732
rect 494848 3720 494854 3732
rect 552658 3720 552664 3732
rect 494848 3692 552664 3720
rect 494848 3680 494854 3692
rect 552658 3680 552664 3692
rect 552716 3680 552722 3732
rect 57422 3612 57428 3664
rect 57480 3652 57486 3664
rect 91554 3652 91560 3664
rect 57480 3624 91560 3652
rect 57480 3612 57486 3624
rect 91554 3612 91560 3624
rect 91612 3612 91618 3664
rect 93946 3612 93952 3664
rect 94004 3652 94010 3664
rect 95142 3652 95148 3664
rect 94004 3624 95148 3652
rect 94004 3612 94010 3624
rect 95142 3612 95148 3624
rect 95200 3612 95206 3664
rect 98638 3612 98644 3664
rect 98696 3652 98702 3664
rect 99282 3652 99288 3664
rect 98696 3624 99288 3652
rect 98696 3612 98702 3624
rect 99282 3612 99288 3624
rect 99340 3612 99346 3664
rect 99834 3612 99840 3664
rect 99892 3652 99898 3664
rect 100662 3652 100668 3664
rect 99892 3624 100668 3652
rect 99892 3612 99898 3624
rect 100662 3612 100668 3624
rect 100720 3612 100726 3664
rect 100757 3655 100815 3661
rect 100757 3621 100769 3655
rect 100803 3652 100815 3655
rect 441798 3652 441804 3664
rect 100803 3624 441804 3652
rect 100803 3621 100815 3624
rect 100757 3615 100815 3621
rect 441798 3612 441804 3624
rect 441856 3612 441862 3664
rect 468478 3612 468484 3664
rect 468536 3652 468542 3664
rect 474550 3652 474556 3664
rect 468536 3624 474556 3652
rect 468536 3612 468542 3624
rect 474550 3612 474556 3624
rect 474608 3612 474614 3664
rect 498838 3612 498844 3664
rect 498896 3652 498902 3664
rect 559742 3652 559748 3664
rect 498896 3624 559748 3652
rect 498896 3612 498902 3624
rect 559742 3612 559748 3624
rect 559800 3612 559806 3664
rect 30098 3544 30104 3596
rect 30156 3584 30162 3596
rect 30156 3556 35894 3584
rect 30156 3544 30162 3556
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3878 3516 3884 3528
rect 2924 3488 3884 3516
rect 2924 3476 2930 3488
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12250 3516 12256 3528
rect 11204 3488 12256 3516
rect 11204 3476 11210 3488
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 26142 3516 26148 3528
rect 25372 3488 26148 3516
rect 25372 3476 25378 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 28902 3516 28908 3528
rect 27764 3488 28908 3516
rect 27764 3476 27770 3488
rect 28902 3476 28908 3488
rect 28960 3476 28966 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 35866 3516 35894 3556
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 37090 3584 37096 3596
rect 36044 3556 37096 3584
rect 36044 3544 36050 3556
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 43070 3544 43076 3596
rect 43128 3584 43134 3596
rect 44082 3584 44088 3596
rect 43128 3556 44088 3584
rect 43128 3544 43134 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45002 3584 45008 3596
rect 44324 3556 45008 3584
rect 44324 3544 44330 3556
rect 45002 3544 45008 3556
rect 45060 3544 45066 3596
rect 55490 3544 55496 3596
rect 55548 3584 55554 3596
rect 56042 3584 56048 3596
rect 55548 3556 56048 3584
rect 55548 3544 55554 3556
rect 56042 3544 56048 3556
rect 56100 3544 56106 3596
rect 59630 3544 59636 3596
rect 59688 3584 59694 3596
rect 78674 3584 78680 3596
rect 59688 3556 78680 3584
rect 59688 3544 59694 3556
rect 78674 3544 78680 3556
rect 78732 3544 78738 3596
rect 82814 3544 82820 3596
rect 82872 3584 82878 3596
rect 83274 3584 83280 3596
rect 82872 3556 83280 3584
rect 82872 3544 82878 3556
rect 83274 3544 83280 3556
rect 83332 3544 83338 3596
rect 84470 3544 84476 3596
rect 84528 3584 84534 3596
rect 442074 3584 442080 3596
rect 84528 3556 442080 3584
rect 84528 3544 84534 3556
rect 442074 3544 442080 3556
rect 442132 3544 442138 3596
rect 456886 3544 456892 3596
rect 456944 3584 456950 3596
rect 458082 3584 458088 3596
rect 456944 3556 458088 3584
rect 456944 3544 456950 3556
rect 458082 3544 458088 3556
rect 458140 3544 458146 3596
rect 473446 3584 473452 3596
rect 470566 3556 473452 3584
rect 394694 3516 394700 3528
rect 35866 3488 394700 3516
rect 394694 3476 394700 3488
rect 394752 3476 394758 3528
rect 396534 3476 396540 3528
rect 396592 3516 396598 3528
rect 397362 3516 397368 3528
rect 396592 3488 397368 3516
rect 396592 3476 396598 3488
rect 397362 3476 397368 3488
rect 397420 3476 397426 3528
rect 398926 3476 398932 3528
rect 398984 3516 398990 3528
rect 399938 3516 399944 3528
rect 398984 3488 399944 3516
rect 398984 3476 398990 3488
rect 399938 3476 399944 3488
rect 399996 3476 400002 3528
rect 403618 3476 403624 3528
rect 403676 3516 403682 3528
rect 404262 3516 404268 3528
rect 403676 3488 404268 3516
rect 403676 3476 403682 3488
rect 404262 3476 404268 3488
rect 404320 3476 404326 3528
rect 406010 3476 406016 3528
rect 406068 3516 406074 3528
rect 407022 3516 407028 3528
rect 406068 3488 407028 3516
rect 406068 3476 406074 3488
rect 407022 3476 407028 3488
rect 407080 3476 407086 3528
rect 408402 3476 408408 3528
rect 408460 3516 408466 3528
rect 441706 3516 441712 3528
rect 408460 3488 441712 3516
rect 408460 3476 408466 3488
rect 441706 3476 441712 3488
rect 441764 3476 441770 3528
rect 448606 3476 448612 3528
rect 448664 3516 448670 3528
rect 449802 3516 449808 3528
rect 448664 3488 449808 3516
rect 448664 3476 448670 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 458818 3476 458824 3528
rect 458876 3516 458882 3528
rect 460382 3516 460388 3528
rect 458876 3488 460388 3516
rect 458876 3476 458882 3488
rect 460382 3476 460388 3488
rect 460440 3476 460446 3528
rect 465718 3476 465724 3528
rect 465776 3516 465782 3528
rect 470566 3516 470594 3556
rect 473446 3544 473452 3556
rect 473504 3544 473510 3596
rect 481634 3544 481640 3596
rect 481692 3584 481698 3596
rect 482830 3584 482836 3596
rect 481692 3556 482836 3584
rect 481692 3544 481698 3556
rect 482830 3544 482836 3556
rect 482888 3544 482894 3596
rect 486510 3544 486516 3596
rect 486568 3584 486574 3596
rect 514754 3584 514760 3596
rect 486568 3556 514760 3584
rect 486568 3544 486574 3556
rect 514754 3544 514760 3556
rect 514812 3544 514818 3596
rect 514864 3556 518894 3584
rect 465776 3488 470594 3516
rect 465776 3476 465782 3488
rect 472710 3476 472716 3528
rect 472768 3516 472774 3528
rect 475746 3516 475752 3528
rect 472768 3488 475752 3516
rect 472768 3476 472774 3488
rect 475746 3476 475752 3488
rect 475804 3476 475810 3528
rect 479518 3476 479524 3528
rect 479576 3516 479582 3528
rect 489914 3516 489920 3528
rect 479576 3488 489920 3516
rect 479576 3476 479582 3488
rect 489914 3476 489920 3488
rect 489972 3476 489978 3528
rect 509878 3476 509884 3528
rect 509936 3516 509942 3528
rect 514864 3516 514892 3556
rect 509936 3488 514892 3516
rect 509936 3476 509942 3488
rect 516778 3476 516784 3528
rect 516836 3516 516842 3528
rect 518342 3516 518348 3528
rect 516836 3488 518348 3516
rect 516836 3476 516842 3488
rect 518342 3476 518348 3488
rect 518400 3476 518406 3528
rect 518866 3516 518894 3556
rect 522298 3544 522304 3596
rect 522356 3584 522362 3596
rect 524230 3584 524236 3596
rect 522356 3556 524236 3584
rect 522356 3544 522362 3556
rect 524230 3544 524236 3556
rect 524288 3544 524294 3596
rect 524325 3587 524383 3593
rect 524325 3553 524337 3587
rect 524371 3584 524383 3587
rect 582190 3584 582196 3596
rect 524371 3556 582196 3584
rect 524371 3553 524383 3556
rect 524325 3547 524383 3553
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 573910 3516 573916 3528
rect 518866 3488 573916 3516
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 14734 3408 14740 3460
rect 14792 3448 14798 3460
rect 397454 3448 397460 3460
rect 14792 3420 397460 3448
rect 14792 3408 14798 3420
rect 397454 3408 397460 3420
rect 397512 3408 397518 3460
rect 404814 3408 404820 3460
rect 404872 3448 404878 3460
rect 441982 3448 441988 3460
rect 404872 3420 441988 3448
rect 404872 3408 404878 3420
rect 441982 3408 441988 3420
rect 442040 3408 442046 3460
rect 461486 3408 461492 3460
rect 461544 3448 461550 3460
rect 495894 3448 495900 3460
rect 461544 3420 495900 3448
rect 461544 3408 461550 3420
rect 495894 3408 495900 3420
rect 495952 3408 495958 3460
rect 507118 3408 507124 3460
rect 507176 3448 507182 3460
rect 570322 3448 570328 3460
rect 507176 3420 570328 3448
rect 507176 3408 507182 3420
rect 570322 3408 570328 3420
rect 570380 3408 570386 3460
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 28960 3352 210648 3380
rect 28960 3340 28966 3352
rect 24210 3272 24216 3324
rect 24268 3312 24274 3324
rect 24268 3284 142154 3312
rect 24268 3272 24274 3284
rect 57238 3204 57244 3256
rect 57296 3244 57302 3256
rect 123478 3244 123484 3256
rect 57296 3216 123484 3244
rect 57296 3204 57302 3216
rect 123478 3204 123484 3216
rect 123536 3204 123542 3256
rect 124674 3204 124680 3256
rect 124732 3244 124738 3256
rect 125502 3244 125508 3256
rect 124732 3216 125508 3244
rect 124732 3204 124738 3216
rect 125502 3204 125508 3216
rect 125560 3204 125566 3256
rect 125870 3204 125876 3256
rect 125928 3244 125934 3256
rect 126790 3244 126796 3256
rect 125928 3216 126796 3244
rect 125928 3204 125934 3216
rect 126790 3204 126796 3216
rect 126848 3204 126854 3256
rect 131758 3204 131764 3256
rect 131816 3244 131822 3256
rect 132402 3244 132408 3256
rect 131816 3216 132408 3244
rect 131816 3204 131822 3216
rect 132402 3204 132408 3216
rect 132460 3204 132466 3256
rect 134150 3204 134156 3256
rect 134208 3244 134214 3256
rect 135162 3244 135168 3256
rect 134208 3216 135168 3244
rect 134208 3204 134214 3216
rect 135162 3204 135168 3216
rect 135220 3204 135226 3256
rect 138842 3204 138848 3256
rect 138900 3244 138906 3256
rect 139302 3244 139308 3256
rect 138900 3216 139308 3244
rect 138900 3204 138906 3216
rect 139302 3204 139308 3216
rect 139360 3204 139366 3256
rect 142126 3244 142154 3284
rect 148318 3272 148324 3324
rect 148376 3312 148382 3324
rect 148962 3312 148968 3324
rect 148376 3284 148968 3312
rect 148376 3272 148382 3284
rect 148962 3272 148968 3284
rect 149020 3272 149026 3324
rect 150618 3272 150624 3324
rect 150676 3312 150682 3324
rect 151722 3312 151728 3324
rect 150676 3284 151728 3312
rect 150676 3272 150682 3284
rect 151722 3272 151728 3284
rect 151780 3272 151786 3324
rect 155402 3272 155408 3324
rect 155460 3312 155466 3324
rect 155862 3312 155868 3324
rect 155460 3284 155868 3312
rect 155460 3272 155466 3284
rect 155862 3272 155868 3284
rect 155920 3272 155926 3324
rect 158898 3272 158904 3324
rect 158956 3312 158962 3324
rect 160002 3312 160008 3324
rect 158956 3284 160008 3312
rect 158956 3272 158962 3284
rect 160002 3272 160008 3284
rect 160060 3272 160066 3324
rect 163682 3272 163688 3324
rect 163740 3312 163746 3324
rect 164142 3312 164148 3324
rect 163740 3284 164148 3312
rect 163740 3272 163746 3284
rect 164142 3272 164148 3284
rect 164200 3272 164206 3324
rect 166074 3272 166080 3324
rect 166132 3312 166138 3324
rect 166902 3312 166908 3324
rect 166132 3284 166908 3312
rect 166132 3272 166138 3284
rect 166902 3272 166908 3284
rect 166960 3272 166966 3324
rect 175458 3272 175464 3324
rect 175516 3312 175522 3324
rect 176562 3312 176568 3324
rect 175516 3284 176568 3312
rect 175516 3272 175522 3284
rect 176562 3272 176568 3284
rect 176620 3272 176626 3324
rect 176654 3272 176660 3324
rect 176712 3312 176718 3324
rect 177850 3312 177856 3324
rect 176712 3284 177856 3312
rect 176712 3272 176718 3284
rect 177850 3272 177856 3284
rect 177908 3272 177914 3324
rect 180242 3272 180248 3324
rect 180300 3312 180306 3324
rect 180702 3312 180708 3324
rect 180300 3284 180708 3312
rect 180300 3272 180306 3284
rect 180702 3272 180708 3284
rect 180760 3272 180766 3324
rect 181438 3272 181444 3324
rect 181496 3312 181502 3324
rect 182082 3312 182088 3324
rect 181496 3284 182088 3312
rect 181496 3272 181502 3284
rect 182082 3272 182088 3284
rect 182140 3272 182146 3324
rect 182542 3272 182548 3324
rect 182600 3312 182606 3324
rect 183462 3312 183468 3324
rect 182600 3284 183468 3312
rect 182600 3272 182606 3284
rect 183462 3272 183468 3284
rect 183520 3272 183526 3324
rect 188522 3272 188528 3324
rect 188580 3312 188586 3324
rect 188982 3312 188988 3324
rect 188580 3284 188988 3312
rect 188580 3272 188586 3284
rect 188982 3272 188988 3284
rect 189040 3272 189046 3324
rect 189718 3272 189724 3324
rect 189776 3312 189782 3324
rect 190362 3312 190368 3324
rect 189776 3284 190368 3312
rect 189776 3272 189782 3284
rect 190362 3272 190368 3284
rect 190420 3272 190426 3324
rect 190822 3272 190828 3324
rect 190880 3312 190886 3324
rect 191742 3312 191748 3324
rect 190880 3284 191748 3312
rect 190880 3272 190886 3284
rect 191742 3272 191748 3284
rect 191800 3272 191806 3324
rect 199102 3272 199108 3324
rect 199160 3312 199166 3324
rect 200022 3312 200028 3324
rect 199160 3284 200028 3312
rect 199160 3272 199166 3284
rect 200022 3272 200028 3284
rect 200080 3272 200086 3324
rect 205082 3272 205088 3324
rect 205140 3312 205146 3324
rect 205542 3312 205548 3324
rect 205140 3284 205548 3312
rect 205140 3272 205146 3284
rect 205542 3272 205548 3284
rect 205600 3272 205606 3324
rect 207382 3272 207388 3324
rect 207440 3312 207446 3324
rect 208210 3312 208216 3324
rect 207440 3284 208216 3312
rect 207440 3272 207446 3284
rect 208210 3272 208216 3284
rect 208268 3272 208274 3324
rect 208578 3272 208584 3324
rect 208636 3312 208642 3324
rect 209682 3312 209688 3324
rect 208636 3284 209688 3312
rect 208636 3272 208642 3284
rect 209682 3272 209688 3284
rect 209740 3272 209746 3324
rect 210620 3312 210648 3352
rect 213362 3340 213368 3392
rect 213420 3380 213426 3392
rect 213822 3380 213828 3392
rect 213420 3352 213828 3380
rect 213420 3340 213426 3352
rect 213822 3340 213828 3352
rect 213880 3340 213886 3392
rect 215662 3340 215668 3392
rect 215720 3380 215726 3392
rect 216582 3380 216588 3392
rect 215720 3352 216588 3380
rect 215720 3340 215726 3352
rect 216582 3340 216588 3352
rect 216640 3340 216646 3392
rect 216858 3340 216864 3392
rect 216916 3380 216922 3392
rect 217962 3380 217968 3392
rect 216916 3352 217968 3380
rect 216916 3340 216922 3352
rect 217962 3340 217968 3352
rect 218020 3340 218026 3392
rect 218054 3340 218060 3392
rect 218112 3380 218118 3392
rect 219342 3380 219348 3392
rect 218112 3352 219348 3380
rect 218112 3340 218118 3352
rect 219342 3340 219348 3352
rect 219400 3340 219406 3392
rect 223942 3340 223948 3392
rect 224000 3380 224006 3392
rect 224678 3380 224684 3392
rect 224000 3352 224684 3380
rect 224000 3340 224006 3352
rect 224678 3340 224684 3352
rect 224736 3340 224742 3392
rect 231026 3340 231032 3392
rect 231084 3380 231090 3392
rect 231762 3380 231768 3392
rect 231084 3352 231768 3380
rect 231084 3340 231090 3352
rect 231762 3340 231768 3352
rect 231820 3340 231826 3392
rect 232222 3340 232228 3392
rect 232280 3380 232286 3392
rect 233142 3380 233148 3392
rect 232280 3352 233148 3380
rect 232280 3340 232286 3352
rect 233142 3340 233148 3352
rect 233200 3340 233206 3392
rect 233418 3340 233424 3392
rect 233476 3380 233482 3392
rect 234522 3380 234528 3392
rect 233476 3352 234528 3380
rect 233476 3340 233482 3352
rect 234522 3340 234528 3352
rect 234580 3340 234586 3392
rect 247586 3340 247592 3392
rect 247644 3380 247650 3392
rect 248322 3380 248328 3392
rect 247644 3352 248328 3380
rect 247644 3340 247650 3352
rect 248322 3340 248328 3352
rect 248380 3340 248386 3392
rect 248782 3340 248788 3392
rect 248840 3380 248846 3392
rect 249702 3380 249708 3392
rect 248840 3352 249708 3380
rect 248840 3340 248846 3352
rect 249702 3340 249708 3352
rect 249760 3340 249766 3392
rect 251174 3340 251180 3392
rect 251232 3380 251238 3392
rect 252462 3380 252468 3392
rect 251232 3352 252468 3380
rect 251232 3340 251238 3352
rect 252462 3340 252468 3352
rect 252520 3340 252526 3392
rect 257062 3340 257068 3392
rect 257120 3380 257126 3392
rect 257982 3380 257988 3392
rect 257120 3352 257988 3380
rect 257120 3340 257126 3352
rect 257982 3340 257988 3352
rect 258040 3340 258046 3392
rect 272426 3340 272432 3392
rect 272484 3380 272490 3392
rect 273162 3380 273168 3392
rect 272484 3352 273168 3380
rect 272484 3340 272490 3352
rect 273162 3340 273168 3352
rect 273220 3340 273226 3392
rect 273622 3340 273628 3392
rect 273680 3380 273686 3392
rect 274542 3380 274548 3392
rect 273680 3352 274548 3380
rect 273680 3340 273686 3352
rect 274542 3340 274548 3352
rect 274600 3340 274606 3392
rect 283098 3340 283104 3392
rect 283156 3380 283162 3392
rect 284202 3380 284208 3392
rect 283156 3352 284208 3380
rect 283156 3340 283162 3352
rect 284202 3340 284208 3352
rect 284260 3340 284266 3392
rect 284294 3340 284300 3392
rect 284352 3380 284358 3392
rect 285582 3380 285588 3392
rect 284352 3352 285588 3380
rect 284352 3340 284358 3352
rect 285582 3340 285588 3352
rect 285640 3340 285646 3392
rect 290182 3340 290188 3392
rect 290240 3380 290246 3392
rect 291102 3380 291108 3392
rect 290240 3352 291108 3380
rect 290240 3340 290246 3352
rect 291102 3340 291108 3352
rect 291160 3340 291166 3392
rect 296070 3340 296076 3392
rect 296128 3380 296134 3392
rect 296622 3380 296628 3392
rect 296128 3352 296628 3380
rect 296128 3340 296134 3352
rect 296622 3340 296628 3352
rect 296680 3340 296686 3392
rect 298462 3340 298468 3392
rect 298520 3380 298526 3392
rect 299382 3380 299388 3392
rect 298520 3352 299388 3380
rect 298520 3340 298526 3352
rect 299382 3340 299388 3352
rect 299440 3340 299446 3392
rect 299474 3340 299480 3392
rect 299532 3380 299538 3392
rect 300762 3380 300768 3392
rect 299532 3352 300768 3380
rect 299532 3340 299538 3352
rect 300762 3340 300768 3352
rect 300820 3340 300826 3392
rect 307757 3383 307815 3389
rect 307757 3349 307769 3383
rect 307803 3380 307815 3383
rect 314654 3380 314660 3392
rect 307803 3352 314660 3380
rect 307803 3349 307815 3352
rect 307757 3343 307815 3349
rect 314654 3340 314660 3352
rect 314712 3340 314718 3392
rect 315022 3340 315028 3392
rect 315080 3380 315086 3392
rect 315942 3380 315948 3392
rect 315080 3352 315948 3380
rect 315080 3340 315086 3352
rect 315942 3340 315948 3352
rect 316000 3340 316006 3392
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 325602 3380 325608 3392
rect 324372 3352 325608 3380
rect 324372 3340 324378 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 331582 3340 331588 3392
rect 331640 3380 331646 3392
rect 332502 3380 332508 3392
rect 331640 3352 332508 3380
rect 331640 3340 331646 3352
rect 332502 3340 332508 3352
rect 332560 3340 332566 3392
rect 345750 3340 345756 3392
rect 345808 3380 345814 3392
rect 346302 3380 346308 3392
rect 345808 3352 346308 3380
rect 345808 3340 345814 3352
rect 346302 3340 346308 3352
rect 346360 3340 346366 3392
rect 354030 3340 354036 3392
rect 354088 3380 354094 3392
rect 354582 3380 354588 3392
rect 354088 3352 354588 3380
rect 354088 3340 354094 3352
rect 354582 3340 354588 3352
rect 354640 3340 354646 3392
rect 357526 3340 357532 3392
rect 357584 3380 357590 3392
rect 358722 3380 358728 3392
rect 357584 3352 358728 3380
rect 357584 3340 357590 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 362310 3340 362316 3392
rect 362368 3380 362374 3392
rect 362862 3380 362868 3392
rect 362368 3352 362868 3380
rect 362368 3340 362374 3352
rect 362862 3340 362868 3352
rect 362920 3340 362926 3392
rect 370590 3340 370596 3392
rect 370648 3380 370654 3392
rect 371142 3380 371148 3392
rect 370648 3352 371148 3380
rect 370648 3340 370654 3352
rect 371142 3340 371148 3352
rect 371200 3340 371206 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 428458 3340 428464 3392
rect 428516 3380 428522 3392
rect 429102 3380 429108 3392
rect 428516 3352 429108 3380
rect 428516 3340 428522 3352
rect 429102 3340 429108 3352
rect 429160 3340 429166 3392
rect 430850 3340 430856 3392
rect 430908 3380 430914 3392
rect 431862 3380 431868 3392
rect 430908 3352 431868 3380
rect 430908 3340 430914 3352
rect 431862 3340 431868 3352
rect 431920 3340 431926 3392
rect 432046 3340 432052 3392
rect 432104 3380 432110 3392
rect 433242 3380 433248 3392
rect 432104 3352 433248 3380
rect 432104 3340 432110 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440234 3340 440240 3392
rect 440292 3380 440298 3392
rect 441522 3380 441528 3392
rect 440292 3352 441528 3380
rect 440292 3340 440298 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 442626 3340 442632 3392
rect 442684 3380 442690 3392
rect 454034 3380 454040 3392
rect 442684 3352 454040 3380
rect 442684 3340 442690 3352
rect 454034 3340 454040 3352
rect 454092 3340 454098 3392
rect 555418 3340 555424 3392
rect 555476 3380 555482 3392
rect 557350 3380 557356 3392
rect 555476 3352 557356 3380
rect 555476 3340 555482 3352
rect 557350 3340 557356 3352
rect 557408 3340 557414 3392
rect 220814 3312 220820 3324
rect 210620 3284 220820 3312
rect 220814 3272 220820 3284
rect 220872 3272 220878 3324
rect 436738 3272 436744 3324
rect 436796 3312 436802 3324
rect 442442 3312 442448 3324
rect 436796 3284 442448 3312
rect 436796 3272 436802 3284
rect 442442 3272 442448 3284
rect 442500 3272 442506 3324
rect 153194 3244 153200 3256
rect 142126 3216 153200 3244
rect 153194 3204 153200 3216
rect 153252 3204 153258 3256
rect 167178 3204 167184 3256
rect 167236 3244 167242 3256
rect 168282 3244 168288 3256
rect 167236 3216 168288 3244
rect 167236 3204 167242 3216
rect 168282 3204 168288 3216
rect 168340 3204 168346 3256
rect 183738 3204 183744 3256
rect 183796 3244 183802 3256
rect 184842 3244 184848 3256
rect 183796 3216 184848 3244
rect 183796 3204 183802 3216
rect 184842 3204 184848 3216
rect 184900 3204 184906 3256
rect 373994 3204 374000 3256
rect 374052 3244 374058 3256
rect 375282 3244 375288 3256
rect 374052 3216 375288 3244
rect 374052 3204 374058 3216
rect 375282 3204 375288 3216
rect 375340 3204 375346 3256
rect 431954 3204 431960 3256
rect 432012 3244 432018 3256
rect 433242 3244 433248 3256
rect 432012 3216 433248 3244
rect 432012 3204 432018 3216
rect 433242 3204 433248 3216
rect 433300 3204 433306 3256
rect 57514 3136 57520 3188
rect 57572 3176 57578 3188
rect 121086 3176 121092 3188
rect 57572 3148 121092 3176
rect 57572 3136 57578 3148
rect 121086 3136 121092 3148
rect 121144 3136 121150 3188
rect 453298 3136 453304 3188
rect 453356 3176 453362 3188
rect 456978 3176 456984 3188
rect 453356 3148 456984 3176
rect 453356 3136 453362 3148
rect 456978 3136 456984 3148
rect 457036 3136 457042 3188
rect 48958 3068 48964 3120
rect 49016 3108 49022 3120
rect 49418 3108 49424 3120
rect 49016 3080 49424 3108
rect 49016 3068 49022 3080
rect 49418 3068 49424 3080
rect 49476 3068 49482 3120
rect 57790 3068 57796 3120
rect 57848 3108 57854 3120
rect 97442 3108 97448 3120
rect 57848 3080 97448 3108
rect 57848 3068 57854 3080
rect 97442 3068 97448 3080
rect 97500 3068 97506 3120
rect 119890 3068 119896 3120
rect 119948 3108 119954 3120
rect 127621 3111 127679 3117
rect 127621 3108 127633 3111
rect 119948 3080 127633 3108
rect 119948 3068 119954 3080
rect 127621 3077 127633 3080
rect 127667 3077 127679 3111
rect 127621 3071 127679 3077
rect 57698 3000 57704 3052
rect 57756 3040 57762 3052
rect 96246 3040 96252 3052
rect 57756 3012 96252 3040
rect 57756 3000 57762 3012
rect 96246 3000 96252 3012
rect 96304 3000 96310 3052
rect 105722 3000 105728 3052
rect 105780 3040 105786 3052
rect 329834 3040 329840 3052
rect 105780 3012 329840 3040
rect 105780 3000 105786 3012
rect 329834 3000 329840 3012
rect 329892 3000 329898 3052
rect 57606 2932 57612 2984
rect 57664 2972 57670 2984
rect 89162 2972 89168 2984
rect 57664 2944 89168 2972
rect 57664 2932 57670 2944
rect 89162 2932 89168 2944
rect 89220 2932 89226 2984
rect 95142 2932 95148 2984
rect 95200 2972 95206 2984
rect 100757 2975 100815 2981
rect 100757 2972 100769 2975
rect 95200 2944 100769 2972
rect 95200 2932 95206 2944
rect 100757 2941 100769 2944
rect 100803 2941 100815 2975
rect 100757 2935 100815 2941
rect 115198 2932 115204 2984
rect 115256 2972 115262 2984
rect 393498 2972 393504 2984
rect 115256 2944 393504 2972
rect 115256 2932 115262 2944
rect 393498 2932 393504 2944
rect 393556 2932 393562 2984
rect 57146 2864 57152 2916
rect 57204 2904 57210 2916
rect 74994 2904 75000 2916
rect 57204 2876 75000 2904
rect 57204 2864 57210 2876
rect 74994 2864 75000 2876
rect 75052 2864 75058 2916
rect 77386 2864 77392 2916
rect 77444 2904 77450 2916
rect 360194 2904 360200 2916
rect 77444 2876 360200 2904
rect 77444 2864 77450 2876
rect 360194 2864 360200 2876
rect 360252 2864 360258 2916
rect 548518 2864 548524 2916
rect 548576 2904 548582 2916
rect 554958 2904 554964 2916
rect 548576 2876 554964 2904
rect 548576 2864 548582 2876
rect 554958 2864 554964 2876
rect 555016 2864 555022 2916
rect 57330 2796 57336 2848
rect 57388 2836 57394 2848
rect 85666 2836 85672 2848
rect 57388 2808 85672 2836
rect 57388 2796 57394 2808
rect 85666 2796 85672 2808
rect 85724 2796 85730 2848
rect 87966 2796 87972 2848
rect 88024 2836 88030 2848
rect 376754 2836 376760 2848
rect 88024 2808 376760 2836
rect 88024 2796 88030 2808
rect 376754 2796 376760 2808
rect 376812 2796 376818 2848
<< via1 >>
rect 144828 700816 144880 700868
rect 170312 700816 170364 700868
rect 92388 700748 92440 700800
rect 202788 700748 202840 700800
rect 57796 700680 57848 700732
rect 154120 700680 154172 700732
rect 172428 700680 172480 700732
rect 300124 700680 300176 700732
rect 122748 700612 122800 700664
rect 235172 700612 235224 700664
rect 283840 700612 283892 700664
rect 439504 700612 439556 700664
rect 137836 700544 137888 700596
rect 305000 700544 305052 700596
rect 429844 700544 429896 700596
rect 440424 700544 440476 700596
rect 57520 700476 57572 700528
rect 332508 700476 332560 700528
rect 348792 700476 348844 700528
rect 439872 700476 439924 700528
rect 464344 700476 464396 700528
rect 478512 700476 478564 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 57612 700408 57664 700460
rect 397460 700408 397512 700460
rect 413652 700408 413704 700460
rect 439780 700408 439832 700460
rect 447784 700408 447836 700460
rect 527180 700408 527232 700460
rect 59268 700340 59320 700392
rect 72976 700340 73028 700392
rect 136548 700340 136600 700392
rect 559656 700340 559708 700392
rect 8116 700272 8168 700324
rect 440608 700272 440660 700324
rect 442356 700272 442408 700324
rect 543464 700272 543516 700324
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 48228 698912 48280 698964
rect 494796 698912 494848 698964
rect 266360 697620 266412 697672
rect 267648 697620 267700 697672
rect 89168 697552 89220 697604
rect 449900 697552 449952 697604
rect 89628 696940 89680 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 440792 683136 440844 683188
rect 3516 670692 3568 670744
rect 439412 670692 439464 670744
rect 442264 670692 442316 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 440332 656888 440384 656940
rect 57704 630640 57756 630692
rect 580172 630640 580224 630692
rect 158628 616836 158680 616888
rect 580172 616836 580224 616888
rect 164148 590656 164200 590708
rect 579620 590656 579672 590708
rect 3516 579640 3568 579692
rect 281540 579640 281592 579692
rect 442448 576852 442500 576904
rect 579620 576852 579672 576904
rect 47952 563048 48004 563100
rect 579896 563048 579948 563100
rect 91560 543532 91612 543584
rect 92388 543532 92440 543584
rect 121828 543532 121880 543584
rect 122748 543532 122800 543584
rect 157892 543532 157944 543584
rect 158628 543532 158680 543584
rect 163044 543532 163096 543584
rect 164148 543532 164200 543584
rect 171416 543532 171468 543584
rect 172428 543532 172480 543584
rect 427084 543328 427136 543380
rect 440516 543328 440568 543380
rect 4068 543260 4120 543312
rect 80612 543260 80664 543312
rect 173992 543260 174044 543312
rect 450084 543260 450136 543312
rect 29644 543192 29696 543244
rect 94780 543192 94832 543244
rect 108304 543192 108356 543244
rect 439596 543192 439648 543244
rect 16488 543124 16540 543176
rect 61292 543124 61344 543176
rect 78036 543124 78088 543176
rect 448612 543124 448664 543176
rect 3700 543056 3752 543108
rect 64512 543056 64564 543108
rect 418712 543056 418764 543108
rect 445852 543056 445904 543108
rect 3516 542988 3568 543040
rect 99932 542988 99984 543040
rect 407764 542988 407816 543040
rect 475384 542988 475436 543040
rect 48136 542920 48188 542972
rect 102508 542920 102560 542972
rect 369768 542920 369820 542972
rect 444380 542920 444432 542972
rect 8208 542852 8260 542904
rect 199108 542852 199160 542904
rect 259644 542852 259696 542904
rect 449992 542852 450044 542904
rect 12348 542784 12400 542836
rect 204260 542784 204312 542836
rect 248696 542784 248748 542836
rect 452660 542784 452712 542836
rect 27528 542716 27580 542768
rect 275744 542716 275796 542768
rect 325332 542716 325384 542768
rect 511264 542716 511316 542768
rect 25504 542648 25556 542700
rect 97356 542648 97408 542700
rect 182364 542648 182416 542700
rect 454132 542648 454184 542700
rect 56692 542580 56744 542632
rect 333704 542580 333756 542632
rect 405188 542580 405240 542632
rect 498844 542580 498896 542632
rect 3240 542512 3292 542564
rect 130200 542512 130252 542564
rect 143724 542512 143776 542564
rect 144828 542512 144880 542564
rect 55036 542444 55088 542496
rect 67088 542444 67140 542496
rect 430304 542444 430356 542496
rect 503720 542444 503772 542496
rect 54300 542376 54352 542428
rect 69664 542376 69716 542428
rect 432880 542376 432932 542428
rect 439688 542376 439740 542428
rect 45376 541628 45428 541680
rect 266360 541628 266412 541680
rect 374920 541560 374972 541612
rect 456984 541560 457036 541612
rect 372344 541492 372396 541544
rect 479524 541492 479576 541544
rect 400036 541424 400088 541476
rect 522304 541424 522356 541476
rect 344652 541356 344704 541408
rect 486424 541356 486476 541408
rect 421932 541288 421984 541340
rect 566464 541288 566516 541340
rect 237748 541220 237800 541272
rect 454040 541220 454092 541272
rect 264796 541152 264848 541204
rect 518164 541152 518216 541204
rect 196532 541084 196584 541136
rect 458824 541084 458876 541136
rect 212632 541016 212684 541068
rect 499580 541016 499632 541068
rect 152096 540948 152148 541000
rect 456800 540948 456852 541000
rect 48044 540268 48096 540320
rect 104900 540268 104952 540320
rect 49516 540200 49568 540252
rect 364340 540200 364392 540252
rect 413560 540175 413612 540184
rect 413560 540141 413569 540175
rect 413569 540141 413603 540175
rect 413603 540141 413612 540175
rect 413560 540132 413612 540141
rect 416136 540175 416188 540184
rect 416136 540141 416145 540175
rect 416145 540141 416179 540175
rect 416179 540141 416188 540175
rect 416136 540132 416188 540141
rect 424508 540175 424560 540184
rect 424508 540141 424517 540175
rect 424517 540141 424551 540175
rect 424551 540141 424560 540175
rect 424508 540132 424560 540141
rect 262220 540107 262272 540116
rect 262220 540073 262229 540107
rect 262229 540073 262263 540107
rect 262263 540073 262272 540107
rect 262220 540064 262272 540073
rect 300860 540107 300912 540116
rect 300860 540073 300869 540107
rect 300869 540073 300903 540107
rect 300903 540073 300912 540107
rect 300860 540064 300912 540073
rect 303436 540107 303488 540116
rect 303436 540073 303445 540107
rect 303445 540073 303479 540107
rect 303479 540073 303488 540107
rect 303436 540064 303488 540073
rect 320180 540107 320232 540116
rect 320180 540073 320189 540107
rect 320189 540073 320223 540107
rect 320223 540073 320232 540107
rect 320180 540064 320232 540073
rect 322756 540107 322808 540116
rect 322756 540073 322765 540107
rect 322765 540073 322799 540107
rect 322799 540073 322808 540107
rect 322756 540064 322808 540073
rect 328552 540107 328604 540116
rect 328552 540073 328561 540107
rect 328561 540073 328595 540107
rect 328595 540073 328604 540107
rect 328552 540064 328604 540073
rect 339500 540107 339552 540116
rect 339500 540073 339509 540107
rect 339509 540073 339543 540107
rect 339543 540073 339552 540107
rect 339500 540064 339552 540073
rect 355600 540107 355652 540116
rect 355600 540073 355609 540107
rect 355609 540073 355643 540107
rect 355643 540073 355652 540107
rect 355600 540064 355652 540073
rect 363972 540064 364024 540116
rect 468484 540064 468536 540116
rect 245384 540039 245436 540048
rect 193680 539928 193732 539980
rect 201960 539971 202012 539980
rect 141424 539860 141476 539912
rect 185952 539835 186004 539844
rect 185952 539801 185961 539835
rect 185961 539801 185995 539835
rect 185995 539801 186004 539835
rect 185952 539792 186004 539801
rect 188528 539835 188580 539844
rect 188528 539801 188537 539835
rect 188537 539801 188571 539835
rect 188571 539801 188580 539835
rect 188528 539792 188580 539801
rect 201960 539937 201969 539971
rect 201969 539937 202003 539971
rect 202003 539937 202012 539971
rect 201960 539928 202012 539937
rect 207204 539971 207256 539980
rect 207204 539937 207213 539971
rect 207213 539937 207247 539971
rect 207247 539937 207256 539971
rect 207204 539928 207256 539937
rect 245384 540005 245393 540039
rect 245393 540005 245427 540039
rect 245427 540005 245436 540039
rect 245384 539996 245436 540005
rect 268384 540039 268436 540048
rect 268384 540005 268393 540039
rect 268393 540005 268427 540039
rect 268427 540005 268436 540039
rect 268384 539996 268436 540005
rect 272892 540039 272944 540048
rect 272892 540005 272901 540039
rect 272901 540005 272935 540039
rect 272935 540005 272944 540039
rect 272892 539996 272944 540005
rect 287152 540039 287204 540048
rect 287152 540005 287161 540039
rect 287161 540005 287195 540039
rect 287195 540005 287204 540039
rect 287152 539996 287204 540005
rect 289820 540039 289872 540048
rect 289820 540005 289829 540039
rect 289829 540005 289863 540039
rect 289863 540005 289872 540039
rect 289820 539996 289872 540005
rect 295248 539996 295300 540048
rect 493324 539996 493376 540048
rect 218704 539971 218756 539980
rect 218704 539937 218713 539971
rect 218713 539937 218747 539971
rect 218747 539937 218756 539971
rect 218704 539928 218756 539937
rect 229744 539971 229796 539980
rect 229744 539937 229753 539971
rect 229753 539937 229787 539971
rect 229787 539937 229796 539971
rect 229744 539928 229796 539937
rect 234436 539928 234488 539980
rect 513380 539928 513432 539980
rect 455420 539860 455472 539912
rect 531412 539792 531464 539844
rect 3332 539724 3384 539776
rect 446036 539724 446088 539776
rect 111248 539656 111300 539708
rect 502340 539656 502392 539708
rect 86776 539588 86828 539640
rect 556252 539588 556304 539640
rect 84016 539563 84068 539572
rect 84016 539529 84025 539563
rect 84025 539529 84059 539563
rect 84059 539529 84068 539563
rect 84016 539520 84068 539529
rect 160744 539520 160796 539572
rect 4804 539452 4856 539504
rect 435180 539452 435232 539504
rect 438400 539520 438452 539572
rect 443000 539520 443052 539572
rect 440240 539452 440292 539504
rect 60648 539384 60700 539436
rect 440976 539384 441028 539436
rect 543740 539316 543792 539368
rect 441068 539248 441120 539300
rect 46848 539180 46900 539232
rect 316960 539180 317012 539232
rect 512000 539180 512052 539232
rect 44088 539112 44140 539164
rect 529940 539112 529992 539164
rect 440884 539044 440936 539096
rect 3516 538976 3568 539028
rect 550640 538976 550692 539028
rect 505100 538908 505152 538960
rect 580172 538840 580224 538892
rect 483020 538772 483072 538824
rect 38568 538704 38620 538756
rect 580540 538704 580592 538756
rect 3884 538636 3936 538688
rect 580908 538636 580960 538688
rect 580724 538568 580776 538620
rect 580632 538500 580684 538552
rect 539692 538432 539744 538484
rect 3700 538364 3752 538416
rect 580080 538364 580132 538416
rect 487160 538296 487212 538348
rect 3976 538228 4028 538280
rect 580448 538228 580500 538280
rect 59820 537888 59872 537940
rect 466460 537888 466512 537940
rect 9588 537820 9640 537872
rect 439964 537820 440016 537872
rect 57336 537752 57388 537804
rect 580908 537752 580960 537804
rect 442080 531292 442132 531344
rect 481640 531292 481692 531344
rect 55128 529932 55180 529984
rect 57428 529932 57480 529984
rect 43996 527144 44048 527196
rect 57336 527144 57388 527196
rect 54944 524424 54996 524476
rect 57336 524424 57388 524476
rect 442540 523608 442592 523660
rect 448520 523608 448572 523660
rect 50988 520276 51040 520328
rect 57336 520276 57388 520328
rect 52368 517488 52420 517540
rect 57336 517488 57388 517540
rect 442908 517488 442960 517540
rect 527824 517488 527876 517540
rect 46756 514768 46808 514820
rect 57336 514768 57388 514820
rect 442908 514768 442960 514820
rect 451280 514768 451332 514820
rect 442908 512184 442960 512236
rect 445944 512184 445996 512236
rect 18604 511980 18656 512032
rect 57336 511980 57388 512032
rect 3424 510552 3476 510604
rect 57152 510552 57204 510604
rect 442540 505112 442592 505164
rect 447140 505112 447192 505164
rect 442816 502324 442868 502376
rect 490012 502324 490064 502376
rect 3332 500964 3384 501016
rect 17224 500964 17276 501016
rect 442540 496816 442592 496868
rect 447508 496816 447560 496868
rect 50896 491308 50948 491360
rect 57612 491308 57664 491360
rect 45468 488520 45520 488572
rect 57612 488520 57664 488572
rect 442724 485800 442776 485852
rect 533344 485800 533396 485852
rect 52092 480224 52144 480276
rect 57612 480224 57664 480276
rect 442908 480224 442960 480276
rect 454684 480224 454736 480276
rect 50804 477504 50856 477556
rect 57060 477504 57112 477556
rect 3424 474716 3476 474768
rect 14464 474716 14516 474768
rect 53748 474716 53800 474768
rect 57612 474716 57664 474768
rect 442908 473356 442960 473408
rect 456892 473356 456944 473408
rect 442908 470568 442960 470620
rect 452752 470568 452804 470620
rect 52000 469208 52052 469260
rect 57612 469208 57664 469260
rect 442908 468664 442960 468716
rect 447600 468664 447652 468716
rect 54852 465060 54904 465112
rect 56876 465060 56928 465112
rect 442816 465060 442868 465112
rect 538864 465060 538916 465112
rect 442908 462544 442960 462596
rect 447232 462544 447284 462596
rect 53656 462340 53708 462392
rect 57612 462340 57664 462392
rect 442908 459824 442960 459876
rect 447416 459824 447468 459876
rect 12256 459552 12308 459604
rect 57612 459552 57664 459604
rect 442908 457104 442960 457156
rect 447324 457104 447376 457156
rect 50712 456764 50764 456816
rect 57612 456764 57664 456816
rect 54668 454044 54720 454096
rect 57612 454044 57664 454096
rect 442908 454044 442960 454096
rect 452844 454044 452896 454096
rect 2688 451256 2740 451308
rect 57612 451256 57664 451308
rect 442908 447448 442960 447500
rect 448704 447448 448756 447500
rect 3976 444388 4028 444440
rect 57060 444388 57112 444440
rect 52276 436092 52328 436144
rect 57612 436092 57664 436144
rect 442724 436092 442776 436144
rect 516784 436092 516836 436144
rect 53564 433304 53616 433356
rect 57612 433304 57664 433356
rect 440976 431876 441028 431928
rect 579988 431876 580040 431928
rect 52184 430584 52236 430636
rect 57612 430584 57664 430636
rect 442908 430584 442960 430636
rect 448796 430584 448848 430636
rect 53380 427796 53432 427848
rect 57612 427796 57664 427848
rect 5448 422288 5500 422340
rect 57612 422288 57664 422340
rect 442908 422288 442960 422340
rect 452936 422288 452988 422340
rect 46664 419500 46716 419552
rect 57612 419500 57664 419552
rect 442540 418888 442592 418940
rect 450176 418888 450228 418940
rect 50620 416780 50672 416832
rect 57612 416780 57664 416832
rect 442724 415624 442776 415676
rect 447692 415624 447744 415676
rect 54760 409844 54812 409896
rect 57520 409844 57572 409896
rect 442540 409844 442592 409896
rect 457076 409844 457128 409896
rect 442540 404608 442592 404660
rect 446128 404608 446180 404660
rect 3608 402908 3660 402960
rect 57520 402908 57572 402960
rect 49608 398828 49660 398880
rect 57520 398828 57572 398880
rect 54208 396040 54260 396092
rect 57520 396040 57572 396092
rect 442908 394952 442960 395004
rect 448888 394952 448940 395004
rect 53472 393320 53524 393372
rect 57520 393320 57572 393372
rect 47860 389172 47912 389224
rect 57520 389172 57572 389224
rect 54484 387812 54536 387864
rect 57520 387812 57572 387864
rect 51908 385024 51960 385076
rect 57520 385024 57572 385076
rect 39304 380876 39356 380928
rect 57520 380876 57572 380928
rect 442908 380876 442960 380928
rect 518900 380876 518952 380928
rect 53104 378156 53156 378208
rect 57520 378156 57572 378208
rect 442908 378156 442960 378208
rect 498200 378156 498252 378208
rect 442908 375368 442960 375420
rect 508504 375368 508556 375420
rect 442908 372784 442960 372836
rect 448980 372784 449032 372836
rect 50528 372580 50580 372632
rect 57520 372580 57572 372632
rect 51540 367072 51592 367124
rect 56876 367072 56928 367124
rect 442908 365712 442960 365764
rect 547880 365712 547932 365764
rect 440884 365644 440936 365696
rect 579988 365644 580040 365696
rect 51816 364352 51868 364404
rect 56876 364352 56928 364404
rect 51724 361564 51776 361616
rect 57520 361564 57572 361616
rect 442632 360544 442684 360596
rect 443644 360544 443696 360596
rect 3792 358708 3844 358760
rect 57520 358708 57572 358760
rect 442724 358368 442776 358420
rect 447876 358368 447928 358420
rect 442908 354696 442960 354748
rect 496820 354696 496872 354748
rect 442908 352384 442960 352436
rect 444564 352384 444616 352436
rect 51632 351908 51684 351960
rect 57520 351908 57572 351960
rect 45284 349120 45336 349172
rect 56876 349120 56928 349172
rect 442724 349120 442776 349172
rect 506572 349120 506624 349172
rect 54024 346400 54076 346452
rect 57520 346400 57572 346452
rect 442908 342592 442960 342644
rect 446312 342592 446364 342644
rect 54576 340892 54628 340944
rect 57520 340892 57572 340944
rect 442908 340892 442960 340944
rect 461584 340892 461636 340944
rect 53288 338104 53340 338156
rect 57520 338104 57572 338156
rect 442908 338104 442960 338156
rect 444656 338104 444708 338156
rect 442724 334160 442776 334212
rect 446220 334160 446272 334212
rect 442908 331576 442960 331628
rect 447968 331576 448020 331628
rect 53196 329808 53248 329860
rect 57520 329808 57572 329860
rect 57520 329196 57572 329248
rect 57888 329196 57940 329248
rect 442908 328448 442960 328500
rect 454224 328448 454276 328500
rect 442540 326068 442592 326120
rect 450268 326068 450320 326120
rect 442540 323076 442592 323128
rect 443552 323076 443604 323128
rect 54392 322940 54444 322992
rect 57336 322940 57388 322992
rect 442908 320152 442960 320204
rect 451372 320152 451424 320204
rect 442908 317500 442960 317552
rect 449072 317500 449124 317552
rect 52828 314644 52880 314696
rect 56876 314644 56928 314696
rect 49424 311856 49476 311908
rect 57336 311856 57388 311908
rect 442724 310768 442776 310820
rect 444472 310768 444524 310820
rect 53012 309136 53064 309188
rect 57336 309136 57388 309188
rect 442908 307776 442960 307828
rect 465724 307776 465776 307828
rect 442448 302472 442500 302524
rect 443276 302472 443328 302524
rect 43904 299480 43956 299532
rect 57336 299480 57388 299532
rect 442908 298052 442960 298104
rect 580908 298052 580960 298104
rect 21364 296692 21416 296744
rect 57336 296692 57388 296744
rect 442448 294584 442500 294636
rect 443368 294584 443420 294636
rect 47768 293972 47820 294024
rect 57888 293972 57940 294024
rect 51264 291184 51316 291236
rect 57060 291184 57112 291236
rect 442908 291184 442960 291236
rect 448060 291184 448112 291236
rect 442908 288464 442960 288516
rect 450360 288464 450412 288516
rect 52736 288396 52788 288448
rect 57336 288396 57388 288448
rect 442908 285744 442960 285796
rect 446404 285744 446456 285796
rect 50436 282888 50488 282940
rect 57336 282888 57388 282940
rect 442816 278740 442868 278792
rect 520924 278740 520976 278792
rect 51448 277380 51500 277432
rect 57336 277380 57388 277432
rect 442540 276632 442592 276684
rect 443460 276632 443512 276684
rect 442908 273232 442960 273284
rect 529204 273232 529256 273284
rect 442908 270784 442960 270836
rect 448244 270784 448296 270836
rect 52644 270512 52696 270564
rect 57336 270512 57388 270564
rect 55680 268064 55732 268116
rect 56600 268064 56652 268116
rect 442908 267724 442960 267776
rect 454316 267724 454368 267776
rect 52920 264936 52972 264988
rect 57428 264936 57480 264988
rect 442908 264936 442960 264988
rect 485044 264936 485096 264988
rect 442908 263168 442960 263220
rect 447784 263168 447836 263220
rect 51356 262216 51408 262268
rect 57428 262216 57480 262268
rect 441068 259360 441120 259412
rect 579804 259360 579856 259412
rect 442908 258068 442960 258120
rect 472624 258068 472676 258120
rect 442540 256504 442592 256556
rect 448152 256504 448204 256556
rect 2780 254056 2832 254108
rect 4896 254056 4948 254108
rect 45192 253920 45244 253972
rect 57428 253920 57480 253972
rect 442908 251132 442960 251184
rect 580816 251132 580868 251184
rect 43812 249772 43864 249824
rect 56876 249772 56928 249824
rect 442724 247052 442776 247104
rect 454408 247052 454460 247104
rect 443644 245556 443696 245608
rect 580172 245556 580224 245608
rect 442908 244264 442960 244316
rect 451556 244264 451608 244316
rect 51172 242904 51224 242956
rect 57336 242904 57388 242956
rect 3056 241408 3108 241460
rect 54300 241408 54352 241460
rect 442724 239096 442776 239148
rect 443828 239096 443880 239148
rect 46572 238756 46624 238808
rect 57336 238756 57388 238808
rect 442908 235968 442960 236020
rect 453028 235968 453080 236020
rect 442908 233384 442960 233436
rect 445760 233384 445812 233436
rect 442908 230664 442960 230716
rect 449164 230664 449216 230716
rect 54300 230460 54352 230512
rect 57336 230460 57388 230512
rect 57336 230324 57388 230376
rect 57888 230324 57940 230376
rect 50344 227740 50396 227792
rect 57888 227740 57940 227792
rect 442908 226312 442960 226364
rect 480260 226312 480312 226364
rect 52552 224952 52604 225004
rect 57888 224952 57940 225004
rect 45100 222164 45152 222216
rect 57888 222164 57940 222216
rect 442632 221008 442684 221060
rect 443644 221008 443696 221060
rect 508504 219376 508556 219428
rect 579988 219376 580040 219428
rect 54116 218016 54168 218068
rect 57888 218016 57940 218068
rect 442908 218016 442960 218068
rect 507860 218016 507912 218068
rect 55772 215296 55824 215348
rect 56600 215296 56652 215348
rect 442908 215296 442960 215348
rect 545764 215296 545816 215348
rect 442724 212848 442776 212900
rect 444012 212848 444064 212900
rect 442724 210264 442776 210316
rect 450452 210264 450504 210316
rect 3516 209788 3568 209840
rect 57888 209788 57940 209840
rect 57796 208496 57848 208548
rect 49516 208292 49568 208344
rect 57704 208292 57756 208344
rect 57796 208292 57848 208344
rect 53932 204280 53984 204332
rect 57704 204280 57756 204332
rect 442908 204212 442960 204264
rect 464344 204212 464396 204264
rect 442908 201492 442960 201544
rect 537484 201492 537536 201544
rect 55588 198704 55640 198756
rect 56600 198704 56652 198756
rect 442908 198704 442960 198756
rect 453120 198704 453172 198756
rect 44916 195984 44968 196036
rect 57704 195984 57756 196036
rect 442908 195304 442960 195356
rect 444748 195304 444800 195356
rect 45376 194488 45428 194540
rect 57704 194488 57756 194540
rect 442908 192584 442960 192636
rect 450544 192584 450596 192636
rect 53840 190476 53892 190528
rect 56876 190476 56928 190528
rect 3332 188980 3384 189032
rect 18604 188980 18656 189032
rect 3240 187620 3292 187672
rect 57704 187620 57756 187672
rect 442632 186464 442684 186516
rect 443736 186464 443788 186516
rect 46480 183540 46532 183592
rect 57704 183540 57756 183592
rect 442908 181024 442960 181076
rect 446496 181024 446548 181076
rect 3976 180820 4028 180872
rect 57704 180820 57756 180872
rect 442908 178304 442960 178356
rect 450636 178304 450688 178356
rect 442724 175584 442776 175636
rect 444840 175584 444892 175636
rect 49516 172524 49568 172576
rect 57704 172524 57756 172576
rect 57796 172456 57848 172508
rect 57796 172252 57848 172304
rect 442908 171096 442960 171148
rect 525800 171096 525852 171148
rect 41328 171028 41380 171080
rect 57888 171028 57940 171080
rect 442908 168376 442960 168428
rect 451648 168376 451700 168428
rect 47676 165588 47728 165640
rect 57888 165588 57940 165640
rect 49332 162868 49384 162920
rect 57888 162868 57940 162920
rect 442908 160624 442960 160676
rect 444932 160624 444984 160676
rect 442724 158652 442776 158704
rect 580816 158652 580868 158704
rect 47952 155864 48004 155916
rect 57888 155864 57940 155916
rect 439504 152464 439556 152516
rect 439596 152464 439648 152516
rect 439504 152260 439556 152312
rect 439596 152260 439648 152312
rect 26148 151784 26200 151836
rect 57888 151784 57940 151836
rect 2780 150084 2832 150136
rect 4804 150084 4856 150136
rect 51080 149200 51132 149252
rect 54208 149200 54260 149252
rect 54208 149064 54260 149116
rect 57888 149064 57940 149116
rect 442908 149064 442960 149116
rect 500960 149064 501012 149116
rect 442816 147568 442868 147620
rect 580908 147568 580960 147620
rect 52460 146616 52512 146668
rect 54024 146616 54076 146668
rect 54024 146276 54076 146328
rect 57888 146276 57940 146328
rect 442908 143624 442960 143676
rect 449256 143624 449308 143676
rect 46296 140768 46348 140820
rect 57888 140768 57940 140820
rect 442908 139408 442960 139460
rect 460204 139408 460256 139460
rect 3332 137912 3384 137964
rect 29644 137912 29696 137964
rect 47952 135260 48004 135312
rect 57888 135260 57940 135312
rect 442908 132064 442960 132116
rect 446588 132064 446640 132116
rect 47584 131112 47636 131164
rect 57888 131112 57940 131164
rect 49240 128324 49292 128376
rect 57888 128324 57940 128376
rect 441528 125604 441580 125656
rect 465080 125604 465132 125656
rect 46388 122816 46440 122868
rect 57888 122816 57940 122868
rect 441528 122816 441580 122868
rect 446772 122816 446824 122868
rect 50252 120096 50304 120148
rect 57888 120096 57940 120148
rect 441528 118668 441580 118720
rect 445024 118668 445076 118720
rect 49148 117308 49200 117360
rect 57888 117308 57940 117360
rect 441528 115948 441580 116000
rect 494704 115948 494756 116000
rect 47492 114520 47544 114572
rect 57888 114520 57940 114572
rect 441528 114384 441580 114436
rect 444104 114384 444156 114436
rect 454684 113092 454736 113144
rect 579988 113092 580040 113144
rect 441528 110440 441580 110492
rect 451464 110440 451516 110492
rect 441528 107652 441580 107704
rect 515404 107652 515456 107704
rect 48228 107584 48280 107636
rect 57888 107584 57940 107636
rect 441528 104864 441580 104916
rect 477500 104864 477552 104916
rect 55496 103504 55548 103556
rect 56600 103504 56652 103556
rect 441528 103436 441580 103488
rect 446036 103436 446088 103488
rect 48044 100648 48096 100700
rect 57888 100648 57940 100700
rect 566464 100648 566516 100700
rect 580172 100648 580224 100700
rect 441528 99356 441580 99408
rect 446680 99356 446732 99408
rect 50160 93848 50212 93900
rect 57888 93848 57940 93900
rect 441528 91060 441580 91112
rect 461676 91060 461728 91112
rect 443920 88000 443972 88052
rect 445024 88000 445076 88052
rect 441528 86980 441580 87032
rect 548524 86980 548576 87032
rect 57888 86003 57940 86012
rect 57888 85969 57897 86003
rect 57897 85969 57931 86003
rect 57931 85969 57940 86003
rect 57888 85960 57940 85969
rect 33048 85552 33100 85604
rect 57888 85552 57940 85604
rect 3332 85484 3384 85536
rect 21364 85484 21416 85536
rect 57888 85459 57940 85468
rect 57888 85425 57897 85459
rect 57897 85425 57931 85459
rect 57931 85425 57940 85459
rect 57888 85416 57940 85425
rect 441528 81404 441580 81456
rect 445024 81404 445076 81456
rect 441528 79976 441580 80028
rect 449900 79976 449952 80028
rect 14464 77188 14516 77240
rect 56876 77188 56928 77240
rect 441528 76304 441580 76356
rect 445116 76304 445168 76356
rect 439504 73176 439556 73228
rect 439504 72972 439556 73024
rect 3516 68416 3568 68468
rect 3700 68416 3752 68468
rect 17224 66172 17276 66224
rect 56876 66172 56928 66224
rect 58072 61752 58124 61804
rect 443552 61752 443604 61804
rect 58992 61684 59044 61736
rect 444012 61684 444064 61736
rect 52092 61616 52144 61668
rect 441252 61616 441304 61668
rect 56324 61548 56376 61600
rect 484400 61548 484452 61600
rect 58440 61480 58492 61532
rect 488540 61480 488592 61532
rect 55588 61412 55640 61464
rect 498292 61412 498344 61464
rect 56232 61344 56284 61396
rect 509240 61344 509292 61396
rect 58624 61276 58676 61328
rect 441160 61276 441212 61328
rect 54024 61208 54076 61260
rect 446312 61208 446364 61260
rect 55680 61140 55732 61192
rect 444104 61140 444156 61192
rect 54484 61072 54536 61124
rect 440516 61072 440568 61124
rect 53840 61004 53892 61056
rect 439688 61004 439740 61056
rect 51540 60936 51592 60988
rect 444656 60936 444708 60988
rect 58532 60868 58584 60920
rect 440792 60868 440844 60920
rect 441528 60868 441580 60920
rect 507124 60868 507176 60920
rect 54668 60800 54720 60852
rect 444840 60800 444892 60852
rect 443184 60732 443236 60784
rect 46664 60664 46716 60716
rect 580540 60664 580592 60716
rect 50252 60596 50304 60648
rect 176660 60596 176712 60648
rect 200028 60596 200080 60648
rect 445944 60596 445996 60648
rect 49608 60528 49660 60580
rect 160100 60528 160152 60580
rect 168288 60528 168340 60580
rect 444564 60528 444616 60580
rect 52000 60460 52052 60512
rect 336740 60460 336792 60512
rect 350448 60503 350500 60512
rect 350448 60469 350457 60503
rect 350457 60469 350491 60503
rect 350491 60469 350500 60503
rect 350448 60460 350500 60469
rect 358728 60460 358780 60512
rect 444932 60460 444984 60512
rect 59912 60392 59964 60444
rect 135260 60392 135312 60444
rect 143540 60435 143592 60444
rect 143540 60401 143549 60435
rect 143549 60401 143583 60435
rect 143583 60401 143592 60435
rect 143540 60392 143592 60401
rect 149152 60435 149204 60444
rect 149152 60401 149161 60435
rect 149161 60401 149195 60435
rect 149195 60401 149204 60435
rect 149152 60392 149204 60401
rect 151728 60392 151780 60444
rect 443828 60392 443880 60444
rect 59268 60324 59320 60376
rect 67640 60324 67692 60376
rect 80060 60367 80112 60376
rect 80060 60333 80069 60367
rect 80069 60333 80103 60367
rect 80103 60333 80112 60367
rect 80060 60324 80112 60333
rect 122748 60324 122800 60376
rect 447968 60324 448020 60376
rect 56692 60256 56744 60308
rect 82820 60256 82872 60308
rect 99288 60256 99340 60308
rect 448244 60256 448296 60308
rect 45008 60188 45060 60240
rect 448152 60188 448204 60240
rect 6828 60120 6880 60172
rect 449072 60120 449124 60172
rect 52644 60052 52696 60104
rect 549260 60052 549312 60104
rect 52828 59984 52880 60036
rect 567200 59984 567252 60036
rect 47584 59916 47636 59968
rect 173900 59916 173952 59968
rect 202788 59916 202840 59968
rect 446404 59916 446456 59968
rect 55956 59848 56008 59900
rect 127164 59848 127216 59900
rect 168380 59891 168432 59900
rect 168380 59857 168389 59891
rect 168389 59857 168423 59891
rect 168423 59857 168432 59891
rect 168380 59848 168432 59857
rect 211068 59891 211120 59900
rect 211068 59857 211077 59891
rect 211077 59857 211111 59891
rect 211111 59857 211120 59891
rect 211068 59848 211120 59857
rect 218060 59891 218112 59900
rect 218060 59857 218069 59891
rect 218069 59857 218103 59891
rect 218103 59857 218112 59891
rect 218060 59848 218112 59857
rect 224684 59891 224736 59900
rect 224684 59857 224693 59891
rect 224693 59857 224727 59891
rect 224727 59857 224736 59891
rect 224684 59848 224736 59857
rect 227628 59848 227680 59900
rect 443000 59848 443052 59900
rect 54852 59780 54904 59832
rect 229192 59780 229244 59832
rect 236000 59823 236052 59832
rect 236000 59789 236009 59823
rect 236009 59789 236043 59823
rect 236043 59789 236052 59823
rect 236000 59780 236052 59789
rect 248328 59780 248380 59832
rect 441344 59780 441396 59832
rect 254032 59755 254084 59764
rect 254032 59721 254041 59755
rect 254041 59721 254075 59755
rect 254075 59721 254084 59755
rect 254032 59712 254084 59721
rect 257988 59755 258040 59764
rect 257988 59721 257997 59755
rect 257997 59721 258031 59755
rect 258031 59721 258040 59755
rect 257988 59712 258040 59721
rect 258080 59755 258132 59764
rect 258080 59721 258089 59755
rect 258089 59721 258123 59755
rect 258123 59721 258132 59755
rect 286968 59755 287020 59764
rect 258080 59712 258132 59721
rect 286968 59721 286977 59755
rect 286977 59721 287011 59755
rect 287011 59721 287020 59755
rect 286968 59712 287020 59721
rect 291108 59755 291160 59764
rect 291108 59721 291117 59755
rect 291117 59721 291151 59755
rect 291151 59721 291160 59755
rect 291108 59712 291160 59721
rect 302240 59755 302292 59764
rect 302240 59721 302249 59755
rect 302249 59721 302283 59755
rect 302283 59721 302292 59755
rect 302240 59712 302292 59721
rect 315948 59755 316000 59764
rect 315948 59721 315957 59755
rect 315957 59721 315991 59755
rect 315991 59721 316000 59755
rect 315948 59712 316000 59721
rect 358820 59755 358872 59764
rect 358820 59721 358829 59755
rect 358829 59721 358863 59755
rect 358863 59721 358872 59755
rect 358820 59712 358872 59721
rect 375380 59755 375432 59764
rect 375380 59721 375389 59755
rect 375389 59721 375423 59755
rect 375423 59721 375432 59755
rect 375380 59712 375432 59721
rect 378048 59755 378100 59764
rect 378048 59721 378057 59755
rect 378057 59721 378091 59755
rect 378091 59721 378100 59755
rect 378048 59712 378100 59721
rect 400128 59755 400180 59764
rect 400128 59721 400137 59755
rect 400137 59721 400171 59755
rect 400171 59721 400180 59755
rect 400128 59712 400180 59721
rect 404268 59755 404320 59764
rect 404268 59721 404277 59755
rect 404277 59721 404311 59755
rect 404311 59721 404320 59755
rect 404268 59712 404320 59721
rect 420920 59712 420972 59764
rect 448612 59712 448664 59764
rect 375288 59687 375340 59696
rect 375288 59653 375297 59687
rect 375297 59653 375331 59687
rect 375331 59653 375340 59687
rect 375288 59644 375340 59653
rect 414020 59644 414072 59696
rect 439596 59644 439648 59696
rect 431868 59619 431920 59628
rect 431868 59585 431877 59619
rect 431877 59585 431911 59619
rect 431911 59585 431920 59619
rect 431868 59576 431920 59585
rect 108948 59372 109000 59424
rect 580172 59372 580224 59424
rect 2964 59304 3016 59356
rect 25504 59304 25556 59356
rect 84476 59304 84528 59356
rect 580448 59304 580500 59356
rect 114744 59236 114796 59288
rect 580264 59236 580316 59288
rect 4896 59168 4948 59220
rect 439320 59168 439372 59220
rect 3792 59100 3844 59152
rect 320824 59100 320876 59152
rect 342720 59100 342772 59152
rect 580632 59100 580684 59152
rect 3608 59032 3660 59084
rect 238392 59032 238444 59084
rect 271236 59032 271288 59084
rect 580816 59032 580868 59084
rect 24768 58964 24820 59016
rect 293132 58964 293184 59016
rect 370412 58964 370464 59016
rect 580356 58964 580408 59016
rect 171048 58896 171100 58948
rect 446128 58896 446180 58948
rect 51264 58828 51316 58880
rect 372620 58828 372672 58880
rect 402888 58828 402940 58880
rect 440700 58828 440752 58880
rect 77208 58760 77260 58812
rect 448060 58760 448112 58812
rect 52736 58692 52788 58744
rect 524420 58692 524472 58744
rect 59084 58624 59136 58676
rect 564532 58624 564584 58676
rect 188988 58556 189040 58608
rect 446496 58556 446548 58608
rect 59728 58488 59780 58540
rect 296720 58488 296772 58540
rect 345940 58488 345992 58540
rect 462320 58488 462372 58540
rect 54208 58420 54260 58472
rect 201500 58420 201552 58472
rect 233148 58420 233200 58472
rect 439412 58420 439464 58472
rect 3884 58352 3936 58404
rect 186228 58352 186280 58404
rect 422300 58352 422352 58404
rect 450084 58352 450136 58404
rect 3516 58284 3568 58336
rect 191380 58284 191432 58336
rect 434720 58284 434772 58336
rect 452660 58284 452712 58336
rect 3424 57876 3476 57928
rect 158536 57876 158588 57928
rect 172704 57876 172756 57928
rect 173808 57876 173860 57928
rect 180432 57876 180484 57928
rect 184940 57876 184992 57928
rect 188804 57876 188856 57928
rect 307760 57876 307812 57928
rect 362868 57876 362920 57928
rect 433524 57876 433576 57928
rect 73528 57808 73580 57860
rect 74448 57808 74500 57860
rect 92848 57808 92900 57860
rect 102232 57808 102284 57860
rect 123116 57808 123168 57860
rect 226524 57808 226576 57860
rect 234528 57808 234580 57860
rect 255136 57808 255188 57860
rect 282184 57808 282236 57860
rect 284208 57808 284260 57860
rect 411628 57808 411680 57860
rect 419540 57808 419592 57860
rect 444380 57808 444432 57860
rect 60004 57740 60056 57792
rect 62580 57672 62632 57724
rect 63316 57672 63368 57724
rect 67732 57672 67784 57724
rect 68928 57672 68980 57724
rect 69756 57740 69808 57792
rect 101220 57740 101272 57792
rect 104808 57740 104860 57792
rect 106372 57740 106424 57792
rect 112168 57740 112220 57792
rect 112996 57740 113048 57792
rect 81532 57672 81584 57724
rect 87052 57672 87104 57724
rect 28908 57604 28960 57656
rect 131488 57740 131540 57792
rect 136640 57740 136692 57792
rect 139216 57604 139268 57656
rect 140044 57604 140096 57656
rect 142436 57740 142488 57792
rect 143448 57740 143500 57792
rect 145012 57740 145064 57792
rect 146208 57740 146260 57792
rect 148968 57740 149020 57792
rect 287980 57740 288032 57792
rect 326620 57740 326672 57792
rect 439044 57740 439096 57792
rect 191840 57672 191892 57724
rect 194600 57672 194652 57724
rect 195888 57672 195940 57724
rect 209872 57672 209924 57724
rect 210700 57672 210752 57724
rect 213828 57672 213880 57724
rect 353668 57672 353720 57724
rect 376208 57672 376260 57724
rect 381544 57672 381596 57724
rect 387156 57672 387208 57724
rect 463700 57672 463752 57724
rect 287060 57604 287112 57656
rect 323400 57604 323452 57656
rect 324228 57604 324280 57656
rect 343548 57604 343600 57656
rect 389732 57604 389784 57656
rect 403256 57604 403308 57656
rect 407764 57604 407816 57656
rect 543004 57604 543056 57656
rect 13728 57536 13780 57588
rect 127900 57536 127952 57588
rect 128268 57536 128320 57588
rect 279608 57536 279660 57588
rect 282184 57536 282236 57588
rect 356888 57536 356940 57588
rect 364340 57536 364392 57588
rect 367836 57536 367888 57588
rect 518256 57536 518308 57588
rect 34428 57468 34480 57520
rect 202972 57468 203024 57520
rect 233240 57468 233292 57520
rect 234436 57468 234488 57520
rect 240968 57468 241020 57520
rect 298744 57468 298796 57520
rect 309876 57468 309928 57520
rect 320824 57468 320876 57520
rect 329196 57468 329248 57520
rect 531964 57468 532016 57520
rect 55036 57400 55088 57452
rect 244280 57400 244332 57452
rect 273168 57400 273220 57452
rect 296352 57400 296404 57452
rect 301504 57400 301556 57452
rect 509884 57400 509936 57452
rect 37188 57332 37240 57384
rect 81900 57332 81952 57384
rect 89628 57332 89680 57384
rect 299480 57332 299532 57384
rect 304724 57332 304776 57384
rect 523684 57332 523736 57384
rect 10968 57264 11020 57316
rect 95424 57264 95476 57316
rect 119896 57264 119948 57316
rect 447784 57264 447836 57316
rect 22008 57196 22060 57248
rect 406476 57196 406528 57248
rect 414204 57196 414256 57248
rect 448612 57196 448664 57248
rect 63408 57128 63460 57180
rect 155960 57128 156012 57180
rect 175280 57128 175332 57180
rect 291200 57128 291252 57180
rect 393228 57128 393280 57180
rect 449256 57128 449308 57180
rect 103796 57060 103848 57112
rect 205640 57060 205692 57112
rect 220728 57060 220780 57112
rect 331772 57060 331824 57112
rect 407028 57060 407080 57112
rect 441068 57060 441120 57112
rect 100668 56992 100720 57044
rect 150164 56992 150216 57044
rect 182088 56992 182140 57044
rect 285404 56992 285456 57044
rect 400680 56992 400732 57044
rect 416780 56992 416832 57044
rect 420000 56992 420052 57044
rect 429200 56992 429252 57044
rect 125692 56924 125744 56976
rect 126888 56924 126940 56976
rect 134064 56924 134116 56976
rect 157340 56924 157392 56976
rect 160008 56924 160060 56976
rect 249340 56924 249392 56976
rect 409052 56924 409104 56976
rect 76104 56856 76156 56908
rect 83464 56856 83516 56908
rect 113088 56856 113140 56908
rect 197176 56856 197228 56908
rect 212448 56856 212500 56908
rect 251916 56856 251968 56908
rect 164148 56788 164200 56840
rect 230020 56788 230072 56840
rect 98000 56720 98052 56772
rect 99196 56720 99248 56772
rect 129648 56720 129700 56772
rect 164332 56720 164384 56772
rect 183652 56720 183704 56772
rect 194692 56720 194744 56772
rect 65156 56652 65208 56704
rect 66076 56652 66128 56704
rect 117320 56584 117372 56636
rect 123484 56584 123536 56636
rect 295984 56584 296036 56636
rect 298928 56584 298980 56636
rect 353208 56516 353260 56568
rect 451280 56516 451332 56568
rect 58164 56448 58216 56500
rect 200120 56448 200172 56500
rect 274548 56448 274600 56500
rect 441436 56448 441488 56500
rect 49240 56380 49292 56432
rect 178040 56380 178092 56432
rect 191748 56380 191800 56432
rect 450636 56380 450688 56432
rect 58256 56312 58308 56364
rect 324320 56312 324372 56364
rect 346308 56312 346360 56364
rect 450452 56312 450504 56364
rect 59820 56244 59872 56296
rect 423680 56244 423732 56296
rect 433248 56244 433300 56296
rect 454224 56244 454276 56296
rect 66168 56176 66220 56228
rect 447600 56176 447652 56228
rect 56968 56108 57020 56160
rect 472716 56108 472768 56160
rect 3424 56040 3476 56092
rect 440056 56040 440108 56092
rect 50160 55972 50212 56024
rect 527180 55972 527232 56024
rect 49516 55904 49568 55956
rect 568580 55904 568632 55956
rect 45468 55836 45520 55888
rect 580264 55836 580316 55888
rect 397368 55768 397420 55820
rect 445116 55768 445168 55820
rect 429108 55700 429160 55752
rect 446680 55700 446732 55752
rect 249708 55020 249760 55072
rect 451556 55020 451608 55072
rect 49148 54952 49200 55004
rect 255320 54952 255372 55004
rect 47952 54884 48004 54936
rect 284300 54884 284352 54936
rect 400036 54884 400088 54936
rect 444748 54884 444800 54936
rect 180708 54816 180760 54868
rect 451372 54816 451424 54868
rect 59636 54748 59688 54800
rect 349160 54748 349212 54800
rect 371148 54748 371200 54800
rect 452936 54748 452988 54800
rect 135168 54680 135220 54732
rect 439964 54680 440016 54732
rect 49332 54612 49384 54664
rect 540980 54612 541032 54664
rect 46756 54544 46808 54596
rect 557540 54544 557592 54596
rect 47768 54476 47820 54528
rect 575480 54476 575532 54528
rect 295248 53524 295300 53576
rect 445024 53524 445076 53576
rect 44916 53456 44968 53508
rect 209780 53456 209832 53508
rect 285588 53456 285640 53508
rect 446588 53456 446640 53508
rect 184848 53388 184900 53440
rect 439780 53388 439832 53440
rect 43996 53320 44048 53372
rect 338120 53320 338172 53372
rect 354588 53320 354640 53372
rect 453120 53320 453172 53372
rect 51172 53252 51224 53304
rect 365720 53252 365772 53304
rect 369768 53252 369820 53304
rect 450544 53252 450596 53304
rect 46480 53184 46532 53236
rect 386420 53184 386472 53236
rect 47492 53116 47544 53168
rect 409880 53116 409932 53168
rect 52552 53048 52604 53100
rect 470600 53048 470652 53100
rect 213920 52028 213972 52080
rect 367100 52028 367152 52080
rect 43904 51960 43956 52012
rect 288440 51960 288492 52012
rect 310428 51960 310480 52012
rect 445852 51960 445904 52012
rect 132408 51892 132460 51944
rect 451648 51892 451700 51944
rect 45100 51824 45152 51876
rect 382280 51824 382332 51876
rect 209872 51756 209924 51808
rect 555424 51756 555476 51808
rect 46296 51688 46348 51740
rect 423772 51688 423824 51740
rect 111708 50532 111760 50584
rect 457076 50532 457128 50584
rect 95148 50464 95200 50516
rect 454408 50464 454460 50516
rect 62028 50396 62080 50448
rect 447508 50396 447560 50448
rect 53380 50328 53432 50380
rect 485780 50328 485832 50380
rect 79968 48968 80020 49020
rect 446772 48968 446824 49020
rect 54944 47540 54996 47592
rect 129740 47540 129792 47592
rect 166908 47540 166960 47592
rect 492680 47540 492732 47592
rect 99196 46860 99248 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 245660 45500 245712 45552
rect 37096 39380 37148 39432
rect 448796 39380 448848 39432
rect 56048 39312 56100 39364
rect 476120 39312 476172 39364
rect 472624 33056 472676 33108
rect 580172 33056 580224 33108
rect 58348 28228 58400 28280
rect 220912 28228 220964 28280
rect 277308 28228 277360 28280
rect 536104 28228 536156 28280
rect 299388 26868 299440 26920
rect 453028 26868 453080 26920
rect 140044 25508 140096 25560
rect 528560 25508 528612 25560
rect 209688 22788 209740 22840
rect 454316 22788 454368 22840
rect 46388 22720 46440 22772
rect 325700 22720 325752 22772
rect 3424 20612 3476 20664
rect 436100 20612 436152 20664
rect 282184 17212 282236 17264
rect 328460 17212 328512 17264
rect 335268 17212 335320 17264
rect 500224 17212 500276 17264
rect 45284 15988 45336 16040
rect 214472 15988 214524 16040
rect 216588 15988 216640 16040
rect 407212 15988 407264 16040
rect 173808 15920 173860 15972
rect 382372 15920 382424 15972
rect 123484 15852 123536 15904
rect 339868 15852 339920 15904
rect 384764 15852 384816 15904
rect 439872 15852 439924 15904
rect 260748 14696 260800 14748
rect 361120 14696 361172 14748
rect 269028 14628 269080 14680
rect 389456 14628 389508 14680
rect 176568 14560 176620 14612
rect 450176 14560 450228 14612
rect 43812 14492 43864 14544
rect 379980 14492 380032 14544
rect 45192 14424 45244 14476
rect 415400 14424 415452 14476
rect 166908 13336 166960 13388
rect 295984 13336 296036 13388
rect 219256 13268 219308 13320
rect 452844 13268 452896 13320
rect 83464 13200 83516 13252
rect 355232 13200 355284 13252
rect 47676 13132 47728 13184
rect 367008 13132 367060 13184
rect 381544 13132 381596 13184
rect 446128 13132 446180 13184
rect 47860 13064 47912 13116
rect 494704 13064 494756 13116
rect 208216 11976 208268 12028
rect 446220 11976 446272 12028
rect 46572 11908 46624 11960
rect 186136 11908 186188 11960
rect 190368 11908 190420 11960
rect 452752 11908 452804 11960
rect 183468 11840 183520 11892
rect 450360 11840 450412 11892
rect 126796 11772 126848 11824
rect 450268 11772 450320 11824
rect 1308 11704 1360 11756
rect 445760 11704 445812 11756
rect 399852 11636 399904 11688
rect 400128 11636 400180 11688
rect 423772 11636 423824 11688
rect 424968 11636 425020 11688
rect 51908 10752 51960 10804
rect 319720 10752 319772 10804
rect 125508 10684 125560 10736
rect 448704 10684 448756 10736
rect 50620 10616 50672 10668
rect 401324 10616 401376 10668
rect 50528 10548 50580 10600
rect 411904 10548 411956 10600
rect 50436 10480 50488 10532
rect 431960 10480 432012 10532
rect 50344 10412 50396 10464
rect 449900 10412 449952 10464
rect 50896 10344 50948 10396
rect 468392 10344 468444 10396
rect 50804 10276 50856 10328
rect 479340 10276 479392 10328
rect 515404 10276 515456 10328
rect 562048 10276 562100 10328
rect 222752 9596 222804 9648
rect 440884 9596 440936 9648
rect 52368 9528 52420 9580
rect 277124 9528 277176 9580
rect 52184 9460 52236 9512
rect 280712 9460 280764 9512
rect 197912 9392 197964 9444
rect 440332 9392 440384 9444
rect 53012 9324 53064 9376
rect 304356 9324 304408 9376
rect 53472 9256 53524 9308
rect 311440 9256 311492 9308
rect 51448 9188 51500 9240
rect 312636 9188 312688 9240
rect 53196 9120 53248 9172
rect 318524 9120 318576 9172
rect 320824 9120 320876 9172
rect 348056 9120 348108 9172
rect 53564 9052 53616 9104
rect 346952 9052 347004 9104
rect 53748 8984 53800 9036
rect 378876 8984 378928 9036
rect 51724 8916 51776 8968
rect 571524 8916 571576 8968
rect 52276 8848 52328 8900
rect 270040 8848 270092 8900
rect 51632 8780 51684 8832
rect 266544 8780 266596 8832
rect 53288 8712 53340 8764
rect 268844 8712 268896 8764
rect 252376 8644 252428 8696
rect 447876 8644 447928 8696
rect 262956 8576 263008 8628
rect 447416 8576 447468 8628
rect 265348 8508 265400 8560
rect 443644 8508 443696 8560
rect 259460 8440 259512 8492
rect 383660 8440 383712 8492
rect 50988 8236 51040 8288
rect 160192 8236 160244 8288
rect 169576 8236 169628 8288
rect 440424 8236 440476 8288
rect 147128 8168 147180 8220
rect 443460 8168 443512 8220
rect 54576 8100 54628 8152
rect 194416 8100 194468 8152
rect 219348 8100 219400 8152
rect 545488 8100 545540 8152
rect 55864 8032 55916 8084
rect 434444 8032 434496 8084
rect 56140 7964 56192 8016
rect 437940 7964 437992 8016
rect 126888 7896 126940 7948
rect 517152 7896 517204 7948
rect 55772 7828 55824 7880
rect 466276 7828 466328 7880
rect 56416 7760 56468 7812
rect 469864 7760 469916 7812
rect 54116 7692 54168 7744
rect 549076 7692 549128 7744
rect 53932 7624 53984 7676
rect 566832 7624 566884 7676
rect 54392 7556 54444 7608
rect 577412 7556 577464 7608
rect 173164 7488 173216 7540
rect 440976 7488 441028 7540
rect 227536 7420 227588 7472
rect 459192 7420 459244 7472
rect 147588 7352 147640 7404
rect 342076 7352 342128 7404
rect 51356 7284 51408 7336
rect 234712 7284 234764 7336
rect 263508 7284 263560 7336
rect 395344 7284 395396 7336
rect 224776 7216 224828 7268
rect 391848 7216 391900 7268
rect 203892 7148 203944 7200
rect 336832 7148 336884 7200
rect 228732 7080 228784 7132
rect 358912 7080 358964 7132
rect 199936 7012 199988 7064
rect 241704 7012 241756 7064
rect 266268 7012 266320 7064
rect 388260 7012 388312 7064
rect 257896 6944 257948 6996
rect 320916 6944 320968 6996
rect 3424 6808 3476 6860
rect 39304 6808 39356 6860
rect 69112 6808 69164 6860
rect 350540 6808 350592 6860
rect 461676 6808 461728 6860
rect 580172 6808 580224 6860
rect 54300 6740 54352 6792
rect 176752 6740 176804 6792
rect 177948 6740 178000 6792
rect 461584 6740 461636 6792
rect 116400 6672 116452 6724
rect 448888 6672 448940 6724
rect 90364 6604 90416 6656
rect 427820 6604 427872 6656
rect 55128 6536 55180 6588
rect 187332 6536 187384 6588
rect 195888 6536 195940 6588
rect 581000 6536 581052 6588
rect 18236 6468 18288 6520
rect 416872 6468 416924 6520
rect 427268 6468 427320 6520
rect 454132 6468 454184 6520
rect 50160 6400 50212 6452
rect 448980 6400 449032 6452
rect 41880 6332 41932 6384
rect 448520 6332 448572 6384
rect 19432 6264 19484 6316
rect 449164 6264 449216 6316
rect 54944 6196 54996 6248
rect 69664 6196 69716 6248
rect 74448 6196 74500 6248
rect 515956 6196 516008 6248
rect 58900 6128 58952 6180
rect 523040 6128 523092 6180
rect 31300 6060 31352 6112
rect 273260 6060 273312 6112
rect 301964 6060 302016 6112
rect 447232 6060 447284 6112
rect 86868 5992 86920 6044
rect 317420 5992 317472 6044
rect 322112 5992 322164 6044
rect 444472 5992 444524 6044
rect 101036 5924 101088 5976
rect 306380 5924 306432 5976
rect 330392 5924 330444 5976
rect 447324 5924 447376 5976
rect 114008 5856 114060 5908
rect 289820 5856 289872 5908
rect 59544 5788 59596 5840
rect 153016 5788 153068 5840
rect 112996 5448 113048 5500
rect 317328 5448 317380 5500
rect 356336 5448 356388 5500
rect 422392 5448 422444 5500
rect 53656 5380 53708 5432
rect 151820 5380 151872 5432
rect 225144 5380 225196 5432
rect 443092 5380 443144 5432
rect 59360 5312 59412 5364
rect 306748 5312 306800 5364
rect 316224 5312 316276 5364
rect 447140 5312 447192 5364
rect 59176 5244 59228 5296
rect 196808 5244 196860 5296
rect 208308 5244 208360 5296
rect 455696 5244 455748 5296
rect 58808 5176 58860 5228
rect 164884 5176 164936 5228
rect 171968 5176 172020 5228
rect 430580 5176 430632 5228
rect 132960 5108 133012 5160
rect 391940 5108 391992 5160
rect 394240 5108 394292 5160
rect 440148 5108 440200 5160
rect 63316 5040 63368 5092
rect 324412 5040 324464 5092
rect 335084 5040 335136 5092
rect 425060 5040 425112 5092
rect 426164 5040 426216 5092
rect 447692 5040 447744 5092
rect 66076 4972 66128 5024
rect 358636 4972 358688 5024
rect 572720 4972 572772 5024
rect 17040 4904 17092 4956
rect 234620 4904 234672 4956
rect 244188 4904 244240 4956
rect 537208 4904 537260 4956
rect 50712 4836 50764 4888
rect 156604 4836 156656 4888
rect 161388 4836 161440 4888
rect 533712 4836 533764 4888
rect 537484 4836 537536 4888
rect 538404 4836 538456 4888
rect 56508 4768 56560 4820
rect 448520 4768 448572 4820
rect 511264 4768 511316 4820
rect 520740 4768 520792 4820
rect 68928 4700 68980 4752
rect 264152 4700 264204 4752
rect 274824 4700 274876 4752
rect 59452 4632 59504 4684
rect 249984 4632 250036 4684
rect 260656 4632 260708 4684
rect 51816 4564 51868 4616
rect 142436 4564 142488 4616
rect 146208 4564 146260 4616
rect 267740 4564 267792 4616
rect 278320 4564 278372 4616
rect 443276 4632 443328 4684
rect 52920 4496 52972 4548
rect 141240 4496 141292 4548
rect 143448 4496 143500 4548
rect 299664 4496 299716 4548
rect 313832 4496 313884 4548
rect 58716 4428 58768 4480
rect 136456 4428 136508 4480
rect 140044 4428 140096 4480
rect 204260 4428 204312 4480
rect 239312 4428 239364 4480
rect 364432 4428 364484 4480
rect 379428 4428 379480 4480
rect 413100 4428 413152 4480
rect 169668 4360 169720 4412
rect 271236 4360 271288 4412
rect 298744 4360 298796 4412
rect 397736 4360 397788 4412
rect 234436 4292 234488 4344
rect 242900 4292 242952 4344
rect 292580 4292 292632 4344
rect 339500 4292 339552 4344
rect 439504 4496 439556 4548
rect 443368 4496 443420 4548
rect 460204 4496 460256 4548
rect 462780 4496 462832 4548
rect 475384 4496 475436 4548
rect 481732 4496 481784 4548
rect 443736 4360 443788 4412
rect 440608 4292 440660 4344
rect 328000 4224 328052 4276
rect 372712 4224 372764 4276
rect 160100 4156 160152 4208
rect 161296 4156 161348 4208
rect 407764 4156 407816 4208
rect 409604 4156 409656 4208
rect 445024 4156 445076 4208
rect 449992 4156 450044 4208
rect 533344 4156 533396 4208
rect 534908 4156 534960 4208
rect 57060 4088 57112 4140
rect 71504 4088 71556 4140
rect 71688 4088 71740 4140
rect 57888 4020 57940 4072
rect 72608 4020 72660 4072
rect 76196 4088 76248 4140
rect 77208 4088 77260 4140
rect 442172 4088 442224 4140
rect 536104 4088 536156 4140
rect 539600 4088 539652 4140
rect 441620 4020 441672 4072
rect 485044 4020 485096 4072
rect 492312 4020 492364 4072
rect 529204 4020 529256 4072
rect 546684 4020 546736 4072
rect 53748 3884 53800 3936
rect 65524 3884 65576 3936
rect 66168 3884 66220 3936
rect 70308 3952 70360 4004
rect 311900 3952 311952 4004
rect 340972 3952 341024 4004
rect 342168 3952 342220 4004
rect 440332 3952 440384 4004
rect 455420 3952 455472 4004
rect 520924 3952 520976 4004
rect 531964 3952 532016 4004
rect 553768 3952 553820 4004
rect 70400 3884 70452 3936
rect 71596 3884 71648 3936
rect 78588 3884 78640 3936
rect 347780 3884 347832 3936
rect 418988 3884 419040 3936
rect 441896 3884 441948 3936
rect 523684 3884 523736 3936
rect 536104 3884 536156 3936
rect 538864 3884 538916 3936
rect 564440 3884 564492 3936
rect 39580 3816 39632 3868
rect 307852 3816 307904 3868
rect 309048 3816 309100 3868
rect 324136 3816 324188 3868
rect 454500 3816 454552 3868
rect 500224 3816 500276 3868
rect 506480 3816 506532 3868
rect 518164 3816 518216 3868
rect 532516 3816 532568 3868
rect 543004 3816 543056 3868
rect 575112 3816 575164 3868
rect 56876 3748 56928 3800
rect 102232 3748 102284 3800
rect 122288 3748 122340 3800
rect 122748 3748 122800 3800
rect 442356 3748 442408 3800
rect 493324 3748 493376 3800
rect 511264 3748 511316 3800
rect 518256 3748 518308 3800
rect 521844 3748 521896 3800
rect 527916 3748 527968 3800
rect 543188 3748 543240 3800
rect 545764 3748 545816 3800
rect 578608 3748 578660 3800
rect 20628 3680 20680 3732
rect 361580 3680 361632 3732
rect 415492 3680 415544 3732
rect 442632 3680 442684 3732
rect 494796 3680 494848 3732
rect 552664 3680 552716 3732
rect 57428 3612 57480 3664
rect 91560 3612 91612 3664
rect 93952 3612 94004 3664
rect 95148 3612 95200 3664
rect 98644 3612 98696 3664
rect 99288 3612 99340 3664
rect 99840 3612 99892 3664
rect 100668 3612 100720 3664
rect 441804 3612 441856 3664
rect 468484 3612 468536 3664
rect 474556 3612 474608 3664
rect 498844 3612 498896 3664
rect 559748 3612 559800 3664
rect 30104 3544 30156 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 2872 3476 2924 3528
rect 3884 3476 3936 3528
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12256 3476 12308 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 25320 3476 25372 3528
rect 26148 3476 26200 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 27712 3476 27764 3528
rect 28908 3476 28960 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 35992 3544 36044 3596
rect 37096 3544 37148 3596
rect 43076 3544 43128 3596
rect 44088 3544 44140 3596
rect 44272 3544 44324 3596
rect 45008 3544 45060 3596
rect 55496 3544 55548 3596
rect 56048 3544 56100 3596
rect 59636 3544 59688 3596
rect 78680 3544 78732 3596
rect 82820 3544 82872 3596
rect 83280 3544 83332 3596
rect 84476 3544 84528 3596
rect 442080 3544 442132 3596
rect 456892 3544 456944 3596
rect 458088 3544 458140 3596
rect 394700 3476 394752 3528
rect 396540 3476 396592 3528
rect 397368 3476 397420 3528
rect 398932 3476 398984 3528
rect 399944 3476 399996 3528
rect 403624 3476 403676 3528
rect 404268 3476 404320 3528
rect 406016 3476 406068 3528
rect 407028 3476 407080 3528
rect 408408 3476 408460 3528
rect 441712 3476 441764 3528
rect 448612 3476 448664 3528
rect 449808 3476 449860 3528
rect 458824 3476 458876 3528
rect 460388 3476 460440 3528
rect 465724 3476 465776 3528
rect 473452 3544 473504 3596
rect 481640 3544 481692 3596
rect 482836 3544 482888 3596
rect 486516 3544 486568 3596
rect 514760 3544 514812 3596
rect 472716 3476 472768 3528
rect 475752 3476 475804 3528
rect 479524 3476 479576 3528
rect 489920 3476 489972 3528
rect 509884 3476 509936 3528
rect 516784 3476 516836 3528
rect 518348 3476 518400 3528
rect 522304 3544 522356 3596
rect 524236 3544 524288 3596
rect 582196 3544 582248 3596
rect 573916 3476 573968 3528
rect 14740 3408 14792 3460
rect 397460 3408 397512 3460
rect 404820 3408 404872 3460
rect 441988 3408 442040 3460
rect 461492 3408 461544 3460
rect 495900 3408 495952 3460
rect 507124 3408 507176 3460
rect 570328 3408 570380 3460
rect 28908 3340 28960 3392
rect 24216 3272 24268 3324
rect 57244 3204 57296 3256
rect 123484 3204 123536 3256
rect 124680 3204 124732 3256
rect 125508 3204 125560 3256
rect 125876 3204 125928 3256
rect 126796 3204 126848 3256
rect 131764 3204 131816 3256
rect 132408 3204 132460 3256
rect 134156 3204 134208 3256
rect 135168 3204 135220 3256
rect 138848 3204 138900 3256
rect 139308 3204 139360 3256
rect 148324 3272 148376 3324
rect 148968 3272 149020 3324
rect 150624 3272 150676 3324
rect 151728 3272 151780 3324
rect 155408 3272 155460 3324
rect 155868 3272 155920 3324
rect 158904 3272 158956 3324
rect 160008 3272 160060 3324
rect 163688 3272 163740 3324
rect 164148 3272 164200 3324
rect 166080 3272 166132 3324
rect 166908 3272 166960 3324
rect 175464 3272 175516 3324
rect 176568 3272 176620 3324
rect 176660 3272 176712 3324
rect 177856 3272 177908 3324
rect 180248 3272 180300 3324
rect 180708 3272 180760 3324
rect 181444 3272 181496 3324
rect 182088 3272 182140 3324
rect 182548 3272 182600 3324
rect 183468 3272 183520 3324
rect 188528 3272 188580 3324
rect 188988 3272 189040 3324
rect 189724 3272 189776 3324
rect 190368 3272 190420 3324
rect 190828 3272 190880 3324
rect 191748 3272 191800 3324
rect 199108 3272 199160 3324
rect 200028 3272 200080 3324
rect 205088 3272 205140 3324
rect 205548 3272 205600 3324
rect 207388 3272 207440 3324
rect 208216 3272 208268 3324
rect 208584 3272 208636 3324
rect 209688 3272 209740 3324
rect 213368 3340 213420 3392
rect 213828 3340 213880 3392
rect 215668 3340 215720 3392
rect 216588 3340 216640 3392
rect 216864 3340 216916 3392
rect 217968 3340 218020 3392
rect 218060 3340 218112 3392
rect 219348 3340 219400 3392
rect 223948 3340 224000 3392
rect 224684 3340 224736 3392
rect 231032 3340 231084 3392
rect 231768 3340 231820 3392
rect 232228 3340 232280 3392
rect 233148 3340 233200 3392
rect 233424 3340 233476 3392
rect 234528 3340 234580 3392
rect 247592 3340 247644 3392
rect 248328 3340 248380 3392
rect 248788 3340 248840 3392
rect 249708 3340 249760 3392
rect 251180 3340 251232 3392
rect 252468 3340 252520 3392
rect 257068 3340 257120 3392
rect 257988 3340 258040 3392
rect 272432 3340 272484 3392
rect 273168 3340 273220 3392
rect 273628 3340 273680 3392
rect 274548 3340 274600 3392
rect 283104 3340 283156 3392
rect 284208 3340 284260 3392
rect 284300 3340 284352 3392
rect 285588 3340 285640 3392
rect 290188 3340 290240 3392
rect 291108 3340 291160 3392
rect 296076 3340 296128 3392
rect 296628 3340 296680 3392
rect 298468 3340 298520 3392
rect 299388 3340 299440 3392
rect 299480 3340 299532 3392
rect 300768 3340 300820 3392
rect 314660 3340 314712 3392
rect 315028 3340 315080 3392
rect 315948 3340 316000 3392
rect 324320 3340 324372 3392
rect 325608 3340 325660 3392
rect 331588 3340 331640 3392
rect 332508 3340 332560 3392
rect 345756 3340 345808 3392
rect 346308 3340 346360 3392
rect 354036 3340 354088 3392
rect 354588 3340 354640 3392
rect 357532 3340 357584 3392
rect 358728 3340 358780 3392
rect 362316 3340 362368 3392
rect 362868 3340 362920 3392
rect 370596 3340 370648 3392
rect 371148 3340 371200 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 428464 3340 428516 3392
rect 429108 3340 429160 3392
rect 430856 3340 430908 3392
rect 431868 3340 431920 3392
rect 432052 3340 432104 3392
rect 433248 3340 433300 3392
rect 440240 3340 440292 3392
rect 441528 3340 441580 3392
rect 442632 3340 442684 3392
rect 454040 3340 454092 3392
rect 555424 3340 555476 3392
rect 557356 3340 557408 3392
rect 220820 3272 220872 3324
rect 436744 3272 436796 3324
rect 442448 3272 442500 3324
rect 153200 3204 153252 3256
rect 167184 3204 167236 3256
rect 168288 3204 168340 3256
rect 183744 3204 183796 3256
rect 184848 3204 184900 3256
rect 374000 3204 374052 3256
rect 375288 3204 375340 3256
rect 431960 3204 432012 3256
rect 433248 3204 433300 3256
rect 57520 3136 57572 3188
rect 121092 3136 121144 3188
rect 453304 3136 453356 3188
rect 456984 3136 457036 3188
rect 48964 3068 49016 3120
rect 49424 3068 49476 3120
rect 57796 3068 57848 3120
rect 97448 3068 97500 3120
rect 119896 3068 119948 3120
rect 57704 3000 57756 3052
rect 96252 3000 96304 3052
rect 105728 3000 105780 3052
rect 329840 3000 329892 3052
rect 57612 2932 57664 2984
rect 89168 2932 89220 2984
rect 95148 2932 95200 2984
rect 115204 2932 115256 2984
rect 393504 2932 393556 2984
rect 57152 2864 57204 2916
rect 75000 2864 75052 2916
rect 77392 2864 77444 2916
rect 360200 2864 360252 2916
rect 548524 2864 548576 2916
rect 554964 2864 555016 2916
rect 57336 2796 57388 2848
rect 85672 2796 85724 2848
rect 87972 2796 88024 2848
rect 376760 2796 376812 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 24320 699718 24348 703520
rect 40512 700466 40540 703520
rect 57796 700732 57848 700738
rect 57796 700674 57848 700680
rect 57520 700528 57572 700534
rect 57520 700470 57572 700476
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3240 542564 3292 542570
rect 3240 542506 3292 542512
rect 3252 527921 3280 542506
rect 3332 539776 3384 539782
rect 3332 539718 3384 539724
rect 3238 527912 3294 527921
rect 3238 527847 3294 527856
rect 3344 514865 3372 539718
rect 3330 514856 3386 514865
rect 3330 514791 3386 514800
rect 3436 510610 3464 632023
rect 3790 619168 3846 619177
rect 3790 619103 3846 619112
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3528 579698 3556 579935
rect 3516 579692 3568 579698
rect 3516 579634 3568 579640
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3528 543046 3556 566879
rect 3516 543040 3568 543046
rect 3516 542982 3568 542988
rect 3516 539028 3568 539034
rect 3516 538970 3568 538976
rect 3424 510604 3476 510610
rect 3424 510546 3476 510552
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 2688 451308 2740 451314
rect 2688 451250 2740 451256
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1320 3534 1348 11698
rect 2700 3534 2728 451250
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 2778 254144 2834 254153
rect 2778 254079 2780 254088
rect 2832 254079 2834 254088
rect 2780 254050 2832 254056
rect 3056 241460 3108 241466
rect 3056 241402 3108 241408
rect 3068 241097 3096 241402
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3146 202872 3202 202881
rect 3146 202807 3202 202816
rect 3160 201929 3188 202807
rect 3146 201920 3202 201929
rect 3146 201855 3202 201864
rect 3344 190454 3372 319223
rect 3252 190426 3372 190454
rect 3252 187678 3280 190426
rect 3332 189032 3384 189038
rect 3332 188974 3384 188980
rect 3344 188873 3372 188974
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3240 187672 3292 187678
rect 3240 187614 3292 187620
rect 2780 150136 2832 150142
rect 2780 150078 2832 150084
rect 2792 149841 2820 150078
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3332 137964 3384 137970
rect 3332 137906 3384 137912
rect 3344 136785 3372 137906
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3146 111752 3202 111761
rect 3146 111687 3202 111696
rect 3160 110673 3188 111687
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 2964 59356 3016 59362
rect 2964 59298 3016 59304
rect 2976 58585 3004 59298
rect 2962 58576 3018 58585
rect 2962 58511 3018 58520
rect 3436 57934 3464 410479
rect 3528 214985 3556 538970
rect 3620 402966 3648 606047
rect 3698 553888 3754 553897
rect 3698 553823 3754 553832
rect 3712 543114 3740 553823
rect 3700 543108 3752 543114
rect 3700 543050 3752 543056
rect 3700 538416 3752 538422
rect 3700 538358 3752 538364
rect 3712 423609 3740 538358
rect 3698 423600 3754 423609
rect 3698 423535 3754 423544
rect 3608 402960 3660 402966
rect 3608 402902 3660 402908
rect 3606 398712 3662 398721
rect 3606 398647 3662 398656
rect 3620 397497 3648 398647
rect 3606 397488 3662 397497
rect 3606 397423 3662 397432
rect 3606 371376 3662 371385
rect 3606 371311 3662 371320
rect 3514 214976 3570 214985
rect 3514 214911 3570 214920
rect 3516 209840 3568 209846
rect 3516 209782 3568 209788
rect 3528 71641 3556 209782
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3516 68468 3568 68474
rect 3516 68410 3568 68416
rect 3528 58342 3556 68410
rect 3620 59090 3648 371311
rect 3804 358766 3832 619103
rect 4068 543312 4120 543318
rect 4068 543254 4120 543260
rect 3884 538688 3936 538694
rect 3884 538630 3936 538636
rect 3792 358760 3844 358766
rect 3792 358702 3844 358708
rect 3698 358456 3754 358465
rect 3698 358391 3754 358400
rect 3712 68474 3740 358391
rect 3790 345400 3846 345409
rect 3790 345335 3846 345344
rect 3700 68468 3752 68474
rect 3700 68410 3752 68416
rect 3804 59158 3832 345335
rect 3896 267209 3924 538630
rect 3976 538280 4028 538286
rect 3976 538222 4028 538228
rect 3988 449585 4016 538222
rect 3974 449576 4030 449585
rect 3974 449511 4030 449520
rect 3976 444440 4028 444446
rect 3976 444382 4028 444388
rect 3988 293185 4016 444382
rect 3974 293176 4030 293185
rect 3974 293111 4030 293120
rect 3882 267200 3938 267209
rect 3882 267135 3938 267144
rect 3976 180872 4028 180878
rect 3976 180814 4028 180820
rect 3882 162888 3938 162897
rect 3882 162823 3938 162832
rect 3792 59152 3844 59158
rect 3792 59094 3844 59100
rect 3608 59084 3660 59090
rect 3608 59026 3660 59032
rect 3896 58410 3924 162823
rect 3884 58404 3936 58410
rect 3884 58346 3936 58352
rect 3516 58336 3568 58342
rect 3516 58278 3568 58284
rect 3424 57928 3476 57934
rect 3424 57870 3476 57876
rect 3424 56092 3476 56098
rect 3424 56034 3476 56040
rect 3436 32473 3464 56034
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3988 6914 4016 180814
rect 3896 6886 4016 6914
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3896 3534 3924 6886
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 584 480 612 3470
rect 1688 480 1716 3470
rect 2884 480 2912 3470
rect 4080 480 4108 543254
rect 16488 543176 16540 543182
rect 16488 543118 16540 543124
rect 8208 542904 8260 542910
rect 8208 542846 8260 542852
rect 4804 539504 4856 539510
rect 4804 539446 4856 539452
rect 4816 150142 4844 539446
rect 5448 422340 5500 422346
rect 5448 422282 5500 422288
rect 4896 254108 4948 254114
rect 4896 254050 4948 254056
rect 4804 150136 4856 150142
rect 4804 150078 4856 150084
rect 4908 59226 4936 254050
rect 4896 59220 4948 59226
rect 4896 59162 4948 59168
rect 5460 6914 5488 422282
rect 6828 60172 6880 60178
rect 6828 60114 6880 60120
rect 6840 6914 6868 60114
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 8220 3534 8248 542846
rect 12348 542836 12400 542842
rect 12348 542778 12400 542784
rect 9588 537872 9640 537878
rect 9588 537814 9640 537820
rect 9600 3534 9628 537814
rect 12256 459604 12308 459610
rect 12256 459546 12308 459552
rect 10968 57316 11020 57322
rect 10968 57258 11020 57264
rect 10980 3534 11008 57258
rect 12268 3534 12296 459546
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 7668 480 7696 3470
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12360 480 12388 542778
rect 14464 474768 14516 474774
rect 14464 474710 14516 474716
rect 14476 77246 14504 474710
rect 14464 77240 14516 77246
rect 14464 77182 14516 77188
rect 13728 57588 13780 57594
rect 13728 57530 13780 57536
rect 13740 6914 13768 57530
rect 13556 6886 13768 6914
rect 13556 480 13584 6886
rect 16500 3534 16528 543118
rect 18604 512032 18656 512038
rect 18604 511974 18656 511980
rect 17224 501016 17276 501022
rect 17224 500958 17276 500964
rect 17236 66230 17264 500958
rect 18616 189038 18644 511974
rect 21364 296744 21416 296750
rect 21364 296686 21416 296692
rect 18604 189032 18656 189038
rect 18604 188974 18656 188980
rect 21376 85542 21404 296686
rect 21364 85536 21416 85542
rect 21364 85478 21416 85484
rect 17224 66224 17276 66230
rect 17224 66166 17276 66172
rect 24780 59022 24808 699654
rect 29644 543244 29696 543250
rect 29644 543186 29696 543192
rect 27528 542768 27580 542774
rect 27528 542710 27580 542716
rect 25504 542700 25556 542706
rect 25504 542642 25556 542648
rect 25516 59362 25544 542642
rect 26148 151836 26200 151842
rect 26148 151778 26200 151784
rect 25504 59356 25556 59362
rect 25504 59298 25556 59304
rect 24768 59016 24820 59022
rect 24768 58958 24820 58964
rect 22008 57248 22060 57254
rect 22008 57190 22060 57196
rect 22020 6914 22048 57190
rect 21836 6886 22048 6914
rect 18236 6520 18288 6526
rect 18236 6462 18288 6468
rect 17040 4956 17092 4962
rect 17040 4898 17092 4904
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14752 480 14780 3402
rect 15948 480 15976 3470
rect 17052 480 17080 4898
rect 18248 480 18276 6462
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19444 480 19472 6258
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20640 480 20668 3674
rect 21836 480 21864 6886
rect 26160 3534 26188 151778
rect 27540 3534 27568 542710
rect 29656 137970 29684 543186
rect 38568 538756 38620 538762
rect 38568 538698 38620 538704
rect 29644 137964 29696 137970
rect 29644 137906 29696 137912
rect 33048 85604 33100 85610
rect 33048 85546 33100 85552
rect 28908 57656 28960 57662
rect 28908 57598 28960 57604
rect 28920 3534 28948 57598
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 30104 3596 30156 3602
rect 30104 3538 30156 3544
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 23018 3360 23074 3369
rect 23018 3295 23074 3304
rect 24216 3324 24268 3330
rect 23032 480 23060 3295
rect 24216 3266 24268 3272
rect 24228 480 24256 3266
rect 25332 480 25360 3470
rect 26528 480 26556 3470
rect 27724 480 27752 3470
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28920 480 28948 3334
rect 30116 480 30144 3538
rect 31312 480 31340 6054
rect 33060 3534 33088 85546
rect 34428 57520 34480 57526
rect 34428 57462 34480 57468
rect 34440 3534 34468 57462
rect 37188 57384 37240 57390
rect 37188 57326 37240 57332
rect 37096 39432 37148 39438
rect 37096 39374 37148 39380
rect 37108 3602 37136 39374
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34794 3496 34850 3505
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34794 3431 34850 3440
rect 34808 480 34836 3431
rect 36004 480 36032 3538
rect 37200 480 37228 57326
rect 38580 6914 38608 538698
rect 39304 380928 39356 380934
rect 39304 380870 39356 380876
rect 38396 6886 38608 6914
rect 38396 480 38424 6886
rect 39316 6866 39344 380870
rect 41340 171086 41368 700402
rect 48228 698964 48280 698970
rect 48228 698906 48280 698912
rect 47952 563100 48004 563106
rect 47952 563042 48004 563048
rect 45376 541680 45428 541686
rect 45376 541622 45428 541628
rect 44088 539164 44140 539170
rect 44088 539106 44140 539112
rect 43996 527196 44048 527202
rect 43996 527138 44048 527144
rect 43904 299532 43956 299538
rect 43904 299474 43956 299480
rect 43812 249824 43864 249830
rect 43812 249766 43864 249772
rect 41328 171080 41380 171086
rect 41328 171022 41380 171028
rect 43824 14550 43852 249766
rect 43916 52018 43944 299474
rect 44008 53378 44036 527138
rect 43996 53372 44048 53378
rect 43996 53314 44048 53320
rect 43904 52012 43956 52018
rect 43904 51954 43956 51960
rect 43812 14544 43864 14550
rect 43812 14486 43864 14492
rect 39304 6860 39356 6866
rect 39304 6802 39356 6808
rect 41880 6384 41932 6390
rect 41880 6326 41932 6332
rect 39580 3868 39632 3874
rect 39580 3810 39632 3816
rect 39592 480 39620 3810
rect 40682 3632 40738 3641
rect 40682 3567 40738 3576
rect 40696 480 40724 3567
rect 41892 480 41920 6326
rect 44100 3602 44128 539106
rect 45284 349172 45336 349178
rect 45284 349114 45336 349120
rect 45192 253972 45244 253978
rect 45192 253914 45244 253920
rect 45100 222216 45152 222222
rect 45100 222158 45152 222164
rect 44916 196036 44968 196042
rect 44916 195978 44968 195984
rect 44928 53514 44956 195978
rect 45008 60240 45060 60246
rect 45008 60182 45060 60188
rect 44916 53508 44968 53514
rect 44916 53450 44968 53456
rect 45020 3602 45048 60182
rect 45112 51882 45140 222158
rect 45100 51876 45152 51882
rect 45100 51818 45152 51824
rect 45204 14482 45232 253914
rect 45296 16046 45324 349114
rect 45388 194546 45416 541622
rect 46848 539232 46900 539238
rect 46848 539174 46900 539180
rect 46756 514820 46808 514826
rect 46756 514762 46808 514768
rect 45468 488572 45520 488578
rect 45468 488514 45520 488520
rect 45376 194540 45428 194546
rect 45376 194482 45428 194488
rect 45480 55894 45508 488514
rect 46664 419552 46716 419558
rect 46664 419494 46716 419500
rect 46572 238808 46624 238814
rect 46572 238750 46624 238756
rect 46480 183592 46532 183598
rect 46480 183534 46532 183540
rect 46296 140820 46348 140826
rect 46296 140762 46348 140768
rect 45468 55888 45520 55894
rect 45468 55830 45520 55836
rect 46308 51746 46336 140762
rect 46388 122868 46440 122874
rect 46388 122810 46440 122816
rect 46296 51740 46348 51746
rect 46296 51682 46348 51688
rect 46400 22778 46428 122810
rect 46492 53242 46520 183534
rect 46480 53236 46532 53242
rect 46480 53178 46532 53184
rect 46388 22772 46440 22778
rect 46388 22714 46440 22720
rect 45284 16040 45336 16046
rect 45284 15982 45336 15988
rect 45192 14476 45244 14482
rect 45192 14418 45244 14424
rect 46584 11966 46612 238750
rect 46676 60722 46704 419494
rect 46664 60716 46716 60722
rect 46664 60658 46716 60664
rect 46768 54602 46796 514762
rect 46756 54596 46808 54602
rect 46756 54538 46808 54544
rect 46572 11960 46624 11966
rect 46572 11902 46624 11908
rect 46860 6914 46888 539174
rect 47860 389224 47912 389230
rect 47860 389166 47912 389172
rect 47768 294024 47820 294030
rect 47768 293966 47820 293972
rect 47676 165640 47728 165646
rect 47676 165582 47728 165588
rect 47584 131164 47636 131170
rect 47584 131106 47636 131112
rect 47492 114572 47544 114578
rect 47492 114514 47544 114520
rect 47504 53174 47532 114514
rect 47596 59974 47624 131106
rect 47584 59968 47636 59974
rect 47584 59910 47636 59916
rect 47492 53168 47544 53174
rect 47492 53110 47544 53116
rect 47688 13190 47716 165582
rect 47780 54534 47808 293966
rect 47768 54528 47820 54534
rect 47768 54470 47820 54476
rect 47676 13184 47728 13190
rect 47676 13126 47728 13132
rect 47872 13122 47900 389166
rect 47964 155922 47992 563042
rect 48136 542972 48188 542978
rect 48136 542914 48188 542920
rect 48044 540320 48096 540326
rect 48044 540262 48096 540268
rect 47952 155916 48004 155922
rect 47952 155858 48004 155864
rect 47952 135312 48004 135318
rect 47952 135254 48004 135260
rect 47964 54942 47992 135254
rect 48056 100706 48084 540262
rect 48044 100700 48096 100706
rect 48044 100642 48096 100648
rect 47952 54936 48004 54942
rect 47952 54878 48004 54884
rect 47860 13116 47912 13122
rect 47860 13058 47912 13064
rect 48148 6914 48176 542914
rect 48240 107642 48268 698906
rect 56692 542632 56744 542638
rect 56692 542574 56744 542580
rect 55036 542496 55088 542502
rect 55036 542438 55088 542444
rect 54300 542428 54352 542434
rect 54300 542370 54352 542376
rect 49516 540252 49568 540258
rect 49516 540194 49568 540200
rect 49424 311908 49476 311914
rect 49424 311850 49476 311856
rect 49332 162920 49384 162926
rect 49332 162862 49384 162868
rect 49240 128376 49292 128382
rect 49240 128318 49292 128324
rect 49148 117360 49200 117366
rect 49148 117302 49200 117308
rect 48228 107636 48280 107642
rect 48228 107578 48280 107584
rect 49160 55010 49188 117302
rect 49252 56438 49280 128318
rect 49240 56432 49292 56438
rect 49240 56374 49292 56380
rect 49148 55004 49200 55010
rect 49148 54946 49200 54952
rect 49344 54670 49372 162862
rect 49332 54664 49384 54670
rect 49332 54606 49384 54612
rect 46676 6886 46888 6914
rect 47872 6886 48176 6914
rect 45466 3768 45522 3777
rect 45466 3703 45522 3712
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 45008 3596 45060 3602
rect 45008 3538 45060 3544
rect 43088 480 43116 3538
rect 44284 480 44312 3538
rect 45480 480 45508 3703
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49436 3126 49464 311850
rect 49528 208350 49556 540194
rect 50988 520328 51040 520334
rect 50988 520270 51040 520276
rect 50896 491360 50948 491366
rect 50896 491302 50948 491308
rect 50804 477556 50856 477562
rect 50804 477498 50856 477504
rect 50712 456816 50764 456822
rect 50712 456758 50764 456764
rect 50620 416832 50672 416838
rect 50620 416774 50672 416780
rect 49608 398880 49660 398886
rect 49608 398822 49660 398828
rect 49516 208344 49568 208350
rect 49516 208286 49568 208292
rect 49516 172576 49568 172582
rect 49516 172518 49568 172524
rect 49528 55962 49556 172518
rect 49620 60586 49648 398822
rect 50528 372632 50580 372638
rect 50528 372574 50580 372580
rect 50436 282940 50488 282946
rect 50436 282882 50488 282888
rect 50344 227792 50396 227798
rect 50344 227734 50396 227740
rect 50252 120148 50304 120154
rect 50252 120090 50304 120096
rect 50160 93900 50212 93906
rect 50160 93842 50212 93848
rect 49608 60580 49660 60586
rect 49608 60522 49660 60528
rect 50172 56030 50200 93842
rect 50264 60654 50292 120090
rect 50252 60648 50304 60654
rect 50252 60590 50304 60596
rect 50160 56024 50212 56030
rect 50160 55966 50212 55972
rect 49516 55956 49568 55962
rect 49516 55898 49568 55904
rect 50356 10470 50384 227734
rect 50448 10538 50476 282882
rect 50540 10606 50568 372574
rect 50632 10674 50660 416774
rect 50620 10668 50672 10674
rect 50620 10610 50672 10616
rect 50528 10600 50580 10606
rect 50528 10542 50580 10548
rect 50436 10532 50488 10538
rect 50436 10474 50488 10480
rect 50344 10464 50396 10470
rect 50344 10406 50396 10412
rect 50160 6452 50212 6458
rect 50160 6394 50212 6400
rect 48964 3120 49016 3126
rect 48964 3062 49016 3068
rect 49424 3120 49476 3126
rect 49424 3062 49476 3068
rect 48976 480 49004 3062
rect 50172 480 50200 6394
rect 50724 4894 50752 456758
rect 50816 10334 50844 477498
rect 50908 10402 50936 491302
rect 50896 10396 50948 10402
rect 50896 10338 50948 10344
rect 50804 10328 50856 10334
rect 50804 10270 50856 10276
rect 51000 8294 51028 520270
rect 52368 517540 52420 517546
rect 52368 517482 52420 517488
rect 52092 480276 52144 480282
rect 52092 480218 52144 480224
rect 52000 469260 52052 469266
rect 52000 469202 52052 469208
rect 51908 385076 51960 385082
rect 51908 385018 51960 385024
rect 51540 367124 51592 367130
rect 51540 367066 51592 367072
rect 51264 291236 51316 291242
rect 51264 291178 51316 291184
rect 51172 242956 51224 242962
rect 51172 242898 51224 242904
rect 51080 149252 51132 149258
rect 51080 149194 51132 149200
rect 50988 8288 51040 8294
rect 50988 8230 51040 8236
rect 51092 6914 51120 149194
rect 51184 53310 51212 242898
rect 51276 58886 51304 291178
rect 51448 277432 51500 277438
rect 51448 277374 51500 277380
rect 51356 262268 51408 262274
rect 51356 262210 51408 262216
rect 51264 58880 51316 58886
rect 51264 58822 51316 58828
rect 51172 53304 51224 53310
rect 51172 53246 51224 53252
rect 51368 7342 51396 262210
rect 51460 9246 51488 277374
rect 51552 60994 51580 367066
rect 51816 364404 51868 364410
rect 51816 364346 51868 364352
rect 51724 361616 51776 361622
rect 51724 361558 51776 361564
rect 51632 351960 51684 351966
rect 51632 351902 51684 351908
rect 51540 60988 51592 60994
rect 51540 60930 51592 60936
rect 51448 9240 51500 9246
rect 51448 9182 51500 9188
rect 51644 8838 51672 351902
rect 51736 8974 51764 361558
rect 51724 8968 51776 8974
rect 51724 8910 51776 8916
rect 51632 8832 51684 8838
rect 51632 8774 51684 8780
rect 51356 7336 51408 7342
rect 51356 7278 51408 7284
rect 51092 6886 51396 6914
rect 50712 4888 50764 4894
rect 50712 4830 50764 4836
rect 51368 480 51396 6886
rect 51828 4622 51856 364346
rect 51920 10810 51948 385018
rect 52012 60518 52040 469202
rect 52104 61674 52132 480218
rect 52276 436144 52328 436150
rect 52276 436086 52328 436092
rect 52184 430636 52236 430642
rect 52184 430578 52236 430584
rect 52092 61668 52144 61674
rect 52092 61610 52144 61616
rect 52000 60512 52052 60518
rect 52000 60454 52052 60460
rect 51908 10804 51960 10810
rect 51908 10746 51960 10752
rect 52196 9518 52224 430578
rect 52184 9512 52236 9518
rect 52184 9454 52236 9460
rect 52288 8906 52316 436086
rect 52380 9586 52408 517482
rect 53748 474768 53800 474774
rect 53748 474710 53800 474716
rect 53656 462392 53708 462398
rect 53656 462334 53708 462340
rect 53564 433356 53616 433362
rect 53564 433298 53616 433304
rect 53380 427848 53432 427854
rect 53380 427790 53432 427796
rect 53104 378208 53156 378214
rect 53104 378150 53156 378156
rect 52828 314696 52880 314702
rect 52828 314638 52880 314644
rect 52736 288448 52788 288454
rect 52736 288390 52788 288396
rect 52644 270564 52696 270570
rect 52644 270506 52696 270512
rect 52552 225004 52604 225010
rect 52552 224946 52604 224952
rect 52460 146668 52512 146674
rect 52460 146610 52512 146616
rect 52472 16574 52500 146610
rect 52564 53106 52592 224946
rect 52656 60110 52684 270506
rect 52644 60104 52696 60110
rect 52644 60046 52696 60052
rect 52748 58750 52776 288390
rect 52840 60042 52868 314638
rect 53012 309188 53064 309194
rect 53012 309130 53064 309136
rect 52920 264988 52972 264994
rect 52920 264930 52972 264936
rect 52828 60036 52880 60042
rect 52828 59978 52880 59984
rect 52736 58744 52788 58750
rect 52736 58686 52788 58692
rect 52552 53100 52604 53106
rect 52552 53042 52604 53048
rect 52472 16546 52592 16574
rect 52368 9580 52420 9586
rect 52368 9522 52420 9528
rect 52276 8900 52328 8906
rect 52276 8842 52328 8848
rect 51816 4616 51868 4622
rect 51816 4558 51868 4564
rect 52564 480 52592 16546
rect 52932 4554 52960 264930
rect 53024 9382 53052 309130
rect 53116 61441 53144 378150
rect 53288 338156 53340 338162
rect 53288 338098 53340 338104
rect 53196 329860 53248 329866
rect 53196 329802 53248 329808
rect 53102 61432 53158 61441
rect 53102 61367 53158 61376
rect 53012 9376 53064 9382
rect 53012 9318 53064 9324
rect 53208 9178 53236 329802
rect 53196 9172 53248 9178
rect 53196 9114 53248 9120
rect 53300 8770 53328 338098
rect 53392 50386 53420 427790
rect 53472 393372 53524 393378
rect 53472 393314 53524 393320
rect 53380 50380 53432 50386
rect 53380 50322 53432 50328
rect 53484 9314 53512 393314
rect 53472 9308 53524 9314
rect 53472 9250 53524 9256
rect 53576 9110 53604 433298
rect 53564 9104 53616 9110
rect 53564 9046 53616 9052
rect 53288 8764 53340 8770
rect 53288 8706 53340 8712
rect 53668 5438 53696 462334
rect 53760 9042 53788 474710
rect 54208 396092 54260 396098
rect 54208 396034 54260 396040
rect 54024 346452 54076 346458
rect 54024 346394 54076 346400
rect 53932 204332 53984 204338
rect 53932 204274 53984 204280
rect 53840 190528 53892 190534
rect 53840 190470 53892 190476
rect 53852 61062 53880 190470
rect 53840 61056 53892 61062
rect 53840 60998 53892 61004
rect 53748 9036 53800 9042
rect 53748 8978 53800 8984
rect 53944 7682 53972 204274
rect 54036 146674 54064 346394
rect 54116 218068 54168 218074
rect 54116 218010 54168 218016
rect 54024 146668 54076 146674
rect 54024 146610 54076 146616
rect 54024 146328 54076 146334
rect 54024 146270 54076 146276
rect 54036 61266 54064 146270
rect 54024 61260 54076 61266
rect 54024 61202 54076 61208
rect 54128 7750 54156 218010
rect 54220 149258 54248 396034
rect 54312 241466 54340 542370
rect 54944 524476 54996 524482
rect 54944 524418 54996 524424
rect 54852 465112 54904 465118
rect 54852 465054 54904 465060
rect 54668 454096 54720 454102
rect 54668 454038 54720 454044
rect 54484 387864 54536 387870
rect 54484 387806 54536 387812
rect 54392 322992 54444 322998
rect 54392 322934 54444 322940
rect 54300 241460 54352 241466
rect 54300 241402 54352 241408
rect 54300 230512 54352 230518
rect 54300 230454 54352 230460
rect 54208 149252 54260 149258
rect 54208 149194 54260 149200
rect 54208 149116 54260 149122
rect 54208 149058 54260 149064
rect 54220 58478 54248 149058
rect 54208 58472 54260 58478
rect 54208 58414 54260 58420
rect 54116 7744 54168 7750
rect 54116 7686 54168 7692
rect 53932 7676 53984 7682
rect 53932 7618 53984 7624
rect 54312 6798 54340 230454
rect 54404 7614 54432 322934
rect 54496 61130 54524 387806
rect 54576 340944 54628 340950
rect 54576 340886 54628 340892
rect 54484 61124 54536 61130
rect 54484 61066 54536 61072
rect 54588 8158 54616 340886
rect 54680 60858 54708 454038
rect 54760 409896 54812 409902
rect 54760 409838 54812 409844
rect 54668 60852 54720 60858
rect 54668 60794 54720 60800
rect 54576 8152 54628 8158
rect 54576 8094 54628 8100
rect 54392 7608 54444 7614
rect 54772 7585 54800 409838
rect 54864 59838 54892 465054
rect 54852 59832 54904 59838
rect 54852 59774 54904 59780
rect 54956 47598 54984 524418
rect 55048 57458 55076 542438
rect 55128 529984 55180 529990
rect 55128 529926 55180 529932
rect 55036 57452 55088 57458
rect 55036 57394 55088 57400
rect 54944 47592 54996 47598
rect 54944 47534 54996 47540
rect 54392 7550 54444 7556
rect 54758 7576 54814 7585
rect 54758 7511 54814 7520
rect 54300 6792 54352 6798
rect 54300 6734 54352 6740
rect 55140 6594 55168 529926
rect 56506 506832 56562 506841
rect 56506 506767 56562 506776
rect 56414 442912 56470 442921
rect 56414 442847 56470 442856
rect 56322 440192 56378 440201
rect 56322 440127 56378 440136
rect 56230 408232 56286 408241
rect 56230 408167 56286 408176
rect 56046 355872 56102 355881
rect 56046 355807 56102 355816
rect 55954 335472 56010 335481
rect 55954 335407 56010 335416
rect 55862 280392 55918 280401
rect 55862 280327 55918 280336
rect 55680 268116 55732 268122
rect 55680 268058 55732 268064
rect 55588 198756 55640 198762
rect 55588 198698 55640 198704
rect 55496 103556 55548 103562
rect 55496 103498 55548 103504
rect 55128 6588 55180 6594
rect 55128 6530 55180 6536
rect 54944 6248 54996 6254
rect 54944 6190 54996 6196
rect 53656 5432 53708 5438
rect 53656 5374 53708 5380
rect 52920 4548 52972 4554
rect 52920 4490 52972 4496
rect 53748 3936 53800 3942
rect 53748 3878 53800 3884
rect 53760 480 53788 3878
rect 54956 480 54984 6190
rect 55508 3602 55536 103498
rect 55600 61470 55628 198698
rect 55588 61464 55640 61470
rect 55588 61406 55640 61412
rect 55692 61198 55720 268058
rect 55772 215348 55824 215354
rect 55772 215290 55824 215296
rect 55680 61192 55732 61198
rect 55680 61134 55732 61140
rect 55784 7886 55812 215290
rect 55876 8090 55904 280327
rect 55968 59906 55996 335407
rect 55956 59900 56008 59906
rect 55956 59842 56008 59848
rect 56060 39370 56088 355807
rect 56138 326632 56194 326641
rect 56138 326567 56194 326576
rect 56048 39364 56100 39370
rect 56048 39306 56100 39312
rect 55864 8084 55916 8090
rect 55864 8026 55916 8032
rect 56152 8022 56180 326567
rect 56244 61402 56272 408167
rect 56336 61606 56364 440127
rect 56324 61600 56376 61606
rect 56324 61542 56376 61548
rect 56232 61396 56284 61402
rect 56232 61338 56284 61344
rect 56140 8016 56192 8022
rect 56140 7958 56192 7964
rect 55772 7880 55824 7886
rect 55772 7822 55824 7828
rect 56428 7818 56456 442847
rect 56416 7812 56468 7818
rect 56416 7754 56468 7760
rect 56520 4826 56548 506767
rect 56598 268832 56654 268841
rect 56598 268767 56654 268776
rect 56612 268122 56640 268767
rect 56600 268116 56652 268122
rect 56600 268058 56652 268064
rect 56598 216472 56654 216481
rect 56598 216407 56654 216416
rect 56612 215354 56640 216407
rect 56600 215348 56652 215354
rect 56600 215290 56652 215296
rect 56598 198792 56654 198801
rect 56598 198727 56600 198736
rect 56652 198727 56654 198736
rect 56600 198698 56652 198704
rect 56598 103592 56654 103601
rect 56598 103527 56600 103536
rect 56652 103527 56654 103536
rect 56600 103498 56652 103504
rect 56704 60314 56732 542574
rect 57336 537804 57388 537810
rect 57336 537746 57388 537752
rect 57348 528554 57376 537746
rect 57428 529984 57480 529990
rect 57426 529952 57428 529961
rect 57480 529952 57482 529961
rect 57426 529887 57482 529896
rect 57348 528526 57468 528554
rect 57334 527232 57390 527241
rect 57334 527167 57336 527176
rect 57388 527167 57390 527176
rect 57336 527138 57388 527144
rect 57334 524512 57390 524521
rect 57334 524447 57336 524456
rect 57388 524447 57390 524456
rect 57336 524418 57388 524424
rect 57334 521112 57390 521121
rect 57334 521047 57390 521056
rect 57348 520334 57376 521047
rect 57336 520328 57388 520334
rect 57336 520270 57388 520276
rect 57334 518392 57390 518401
rect 57334 518327 57390 518336
rect 57348 517546 57376 518327
rect 57336 517540 57388 517546
rect 57336 517482 57388 517488
rect 57334 515672 57390 515681
rect 57334 515607 57390 515616
rect 57348 514826 57376 515607
rect 57336 514820 57388 514826
rect 57336 514762 57388 514768
rect 57334 512952 57390 512961
rect 57334 512887 57390 512896
rect 57348 512038 57376 512887
rect 57336 512032 57388 512038
rect 57336 511974 57388 511980
rect 57152 510604 57204 510610
rect 57152 510546 57204 510552
rect 57164 509561 57192 510546
rect 57150 509552 57206 509561
rect 57150 509487 57206 509496
rect 57058 477592 57114 477601
rect 57058 477527 57060 477536
rect 57112 477527 57114 477536
rect 57060 477498 57112 477504
rect 56874 466032 56930 466041
rect 56874 465967 56930 465976
rect 56888 465118 56916 465967
rect 56876 465112 56928 465118
rect 56876 465054 56928 465060
rect 57058 445632 57114 445641
rect 57058 445567 57114 445576
rect 57072 444446 57100 445567
rect 57060 444440 57112 444446
rect 57060 444382 57112 444388
rect 56874 367432 56930 367441
rect 56874 367367 56930 367376
rect 56888 367130 56916 367367
rect 56876 367124 56928 367130
rect 56876 367066 56928 367072
rect 56874 364712 56930 364721
rect 56874 364647 56930 364656
rect 56888 364410 56916 364647
rect 56876 364404 56928 364410
rect 56876 364346 56928 364352
rect 56874 350432 56930 350441
rect 56874 350367 56930 350376
rect 56888 349178 56916 350367
rect 56876 349172 56928 349178
rect 56876 349114 56928 349120
rect 57334 323912 57390 323921
rect 57334 323847 57390 323856
rect 57348 322998 57376 323847
rect 57336 322992 57388 322998
rect 57336 322934 57388 322940
rect 56874 315072 56930 315081
rect 56874 315007 56930 315016
rect 56888 314702 56916 315007
rect 56876 314696 56928 314702
rect 56876 314638 56928 314644
rect 57334 312352 57390 312361
rect 57334 312287 57390 312296
rect 57348 311914 57376 312287
rect 57336 311908 57388 311914
rect 57336 311850 57388 311856
rect 57334 309632 57390 309641
rect 57334 309567 57390 309576
rect 57348 309194 57376 309567
rect 57336 309188 57388 309194
rect 57336 309130 57388 309136
rect 57334 300792 57390 300801
rect 57334 300727 57390 300736
rect 57348 299538 57376 300727
rect 57336 299532 57388 299538
rect 57336 299474 57388 299480
rect 57334 298072 57390 298081
rect 57334 298007 57390 298016
rect 57348 296750 57376 298007
rect 57336 296744 57388 296750
rect 57336 296686 57388 296692
rect 57058 291952 57114 291961
rect 57058 291887 57114 291896
rect 57072 291242 57100 291887
rect 57060 291236 57112 291242
rect 57060 291178 57112 291184
rect 57334 289232 57390 289241
rect 57334 289167 57390 289176
rect 57348 288454 57376 289167
rect 57336 288448 57388 288454
rect 57336 288390 57388 288396
rect 57334 283112 57390 283121
rect 57334 283047 57390 283056
rect 57348 282946 57376 283047
rect 57336 282940 57388 282946
rect 57336 282882 57388 282888
rect 57334 277672 57390 277681
rect 57334 277607 57390 277616
rect 57348 277438 57376 277607
rect 57336 277432 57388 277438
rect 57336 277374 57388 277380
rect 57334 271552 57390 271561
rect 57334 271487 57390 271496
rect 57348 270570 57376 271487
rect 57336 270564 57388 270570
rect 57336 270506 57388 270512
rect 57440 267734 57468 528526
rect 57532 504121 57560 700470
rect 57612 700460 57664 700466
rect 57612 700402 57664 700408
rect 57518 504112 57574 504121
rect 57518 504047 57574 504056
rect 57624 495281 57652 700402
rect 57704 630692 57756 630698
rect 57704 630634 57756 630640
rect 57610 495272 57666 495281
rect 57610 495207 57666 495216
rect 57610 492552 57666 492561
rect 57610 492487 57666 492496
rect 57624 491366 57652 492487
rect 57612 491360 57664 491366
rect 57612 491302 57664 491308
rect 57610 489152 57666 489161
rect 57610 489087 57666 489096
rect 57624 488578 57652 489087
rect 57612 488572 57664 488578
rect 57612 488514 57664 488520
rect 57610 480992 57666 481001
rect 57610 480927 57666 480936
rect 57624 480282 57652 480927
rect 57612 480276 57664 480282
rect 57612 480218 57664 480224
rect 57610 474872 57666 474881
rect 57610 474807 57666 474816
rect 57624 474774 57652 474807
rect 57612 474768 57664 474774
rect 57612 474710 57664 474716
rect 57610 469432 57666 469441
rect 57610 469367 57666 469376
rect 57624 469266 57652 469367
rect 57612 469260 57664 469266
rect 57612 469202 57664 469208
rect 57610 463312 57666 463321
rect 57610 463247 57666 463256
rect 57624 462398 57652 463247
rect 57612 462392 57664 462398
rect 57612 462334 57664 462340
rect 57610 460592 57666 460601
rect 57610 460527 57666 460536
rect 57624 459610 57652 460527
rect 57612 459604 57664 459610
rect 57612 459546 57664 459552
rect 57610 457872 57666 457881
rect 57610 457807 57666 457816
rect 57624 456822 57652 457807
rect 57612 456816 57664 456822
rect 57612 456758 57664 456764
rect 57610 454472 57666 454481
rect 57610 454407 57666 454416
rect 57624 454102 57652 454407
rect 57612 454096 57664 454102
rect 57612 454038 57664 454044
rect 57610 451752 57666 451761
rect 57610 451687 57666 451696
rect 57624 451314 57652 451687
rect 57612 451308 57664 451314
rect 57612 451250 57664 451256
rect 57610 437472 57666 437481
rect 57610 437407 57666 437416
rect 57624 436150 57652 437407
rect 57612 436144 57664 436150
rect 57612 436086 57664 436092
rect 57610 434072 57666 434081
rect 57610 434007 57666 434016
rect 57624 433362 57652 434007
rect 57612 433356 57664 433362
rect 57612 433298 57664 433304
rect 57610 431352 57666 431361
rect 57610 431287 57666 431296
rect 57624 430642 57652 431287
rect 57612 430636 57664 430642
rect 57612 430578 57664 430584
rect 57610 428632 57666 428641
rect 57610 428567 57666 428576
rect 57624 427854 57652 428567
rect 57612 427848 57664 427854
rect 57612 427790 57664 427796
rect 57610 422512 57666 422521
rect 57610 422447 57666 422456
rect 57624 422346 57652 422447
rect 57612 422340 57664 422346
rect 57612 422282 57664 422288
rect 57610 419792 57666 419801
rect 57610 419727 57666 419736
rect 57624 419558 57652 419727
rect 57612 419552 57664 419558
rect 57612 419494 57664 419500
rect 57610 417072 57666 417081
rect 57610 417007 57666 417016
rect 57624 416838 57652 417007
rect 57612 416832 57664 416838
rect 57612 416774 57664 416780
rect 57610 413672 57666 413681
rect 57610 413607 57666 413616
rect 57518 410952 57574 410961
rect 57518 410887 57574 410896
rect 57532 409902 57560 410887
rect 57520 409896 57572 409902
rect 57520 409838 57572 409844
rect 57520 402960 57572 402966
rect 57520 402902 57572 402908
rect 57532 402121 57560 402902
rect 57518 402112 57574 402121
rect 57518 402047 57574 402056
rect 57518 399392 57574 399401
rect 57518 399327 57574 399336
rect 57532 398886 57560 399327
rect 57520 398880 57572 398886
rect 57520 398822 57572 398828
rect 57518 396672 57574 396681
rect 57518 396607 57574 396616
rect 57532 396098 57560 396607
rect 57520 396092 57572 396098
rect 57520 396034 57572 396040
rect 57518 393952 57574 393961
rect 57518 393887 57574 393896
rect 57532 393378 57560 393887
rect 57520 393372 57572 393378
rect 57520 393314 57572 393320
rect 57518 390552 57574 390561
rect 57518 390487 57574 390496
rect 57532 389230 57560 390487
rect 57520 389224 57572 389230
rect 57520 389166 57572 389172
rect 57520 387864 57572 387870
rect 57518 387832 57520 387841
rect 57572 387832 57574 387841
rect 57518 387767 57574 387776
rect 57518 385112 57574 385121
rect 57518 385047 57520 385056
rect 57572 385047 57574 385056
rect 57520 385018 57572 385024
rect 57518 381712 57574 381721
rect 57518 381647 57574 381656
rect 57532 380934 57560 381647
rect 57520 380928 57572 380934
rect 57520 380870 57572 380876
rect 57518 378992 57574 379001
rect 57518 378927 57574 378936
rect 57532 378214 57560 378927
rect 57520 378208 57572 378214
rect 57520 378150 57572 378156
rect 57518 373552 57574 373561
rect 57518 373487 57574 373496
rect 57532 372638 57560 373487
rect 57520 372632 57572 372638
rect 57520 372574 57572 372580
rect 57518 361992 57574 362001
rect 57518 361927 57574 361936
rect 57532 361622 57560 361927
rect 57520 361616 57572 361622
rect 57520 361558 57572 361564
rect 57520 358760 57572 358766
rect 57520 358702 57572 358708
rect 57532 358601 57560 358702
rect 57518 358592 57574 358601
rect 57518 358527 57574 358536
rect 57518 353152 57574 353161
rect 57518 353087 57574 353096
rect 57532 351966 57560 353087
rect 57520 351960 57572 351966
rect 57520 351902 57572 351908
rect 57518 347032 57574 347041
rect 57518 346967 57574 346976
rect 57532 346458 57560 346967
rect 57520 346452 57572 346458
rect 57520 346394 57572 346400
rect 57518 341592 57574 341601
rect 57518 341527 57574 341536
rect 57532 340950 57560 341527
rect 57520 340944 57572 340950
rect 57520 340886 57572 340892
rect 57518 338192 57574 338201
rect 57518 338127 57520 338136
rect 57572 338127 57574 338136
rect 57520 338098 57572 338104
rect 57518 330032 57574 330041
rect 57518 329967 57574 329976
rect 57532 329866 57560 329967
rect 57520 329860 57572 329866
rect 57520 329802 57572 329808
rect 57520 329248 57572 329254
rect 57520 329190 57572 329196
rect 57348 267706 57468 267734
rect 57348 260001 57376 267706
rect 57426 266112 57482 266121
rect 57426 266047 57482 266056
rect 57440 264994 57468 266047
rect 57428 264988 57480 264994
rect 57428 264930 57480 264936
rect 57426 262712 57482 262721
rect 57426 262647 57482 262656
rect 57440 262274 57468 262647
rect 57428 262268 57480 262274
rect 57428 262210 57480 262216
rect 57334 259992 57390 260001
rect 57334 259927 57390 259936
rect 57426 254552 57482 254561
rect 57426 254487 57482 254496
rect 57440 253978 57468 254487
rect 57428 253972 57480 253978
rect 57428 253914 57480 253920
rect 56874 251152 56930 251161
rect 56874 251087 56930 251096
rect 56888 249830 56916 251087
rect 56876 249824 56928 249830
rect 56876 249766 56928 249772
rect 57426 248432 57482 248441
rect 57426 248367 57482 248376
rect 57334 242992 57390 243001
rect 57334 242927 57336 242936
rect 57388 242927 57390 242936
rect 57336 242898 57388 242904
rect 57334 239592 57390 239601
rect 57334 239527 57390 239536
rect 57348 238814 57376 239527
rect 57336 238808 57388 238814
rect 57336 238750 57388 238756
rect 57242 234152 57298 234161
rect 57242 234087 57298 234096
rect 56874 190632 56930 190641
rect 56874 190567 56930 190576
rect 56888 190534 56916 190567
rect 56876 190528 56928 190534
rect 56876 190470 56928 190476
rect 57150 158672 57206 158681
rect 57150 158607 57206 158616
rect 57058 143712 57114 143721
rect 57058 143647 57114 143656
rect 56966 126712 57022 126721
rect 56966 126647 57022 126656
rect 56876 77240 56928 77246
rect 56876 77182 56928 77188
rect 56888 77081 56916 77182
rect 56874 77072 56930 77081
rect 56874 77007 56930 77016
rect 56782 71632 56838 71641
rect 56782 71567 56838 71576
rect 56796 64874 56824 71567
rect 56876 66224 56928 66230
rect 56876 66166 56928 66172
rect 56888 65521 56916 66166
rect 56874 65512 56930 65521
rect 56874 65447 56930 65456
rect 56796 64846 56916 64874
rect 56692 60308 56744 60314
rect 56692 60250 56744 60256
rect 56508 4820 56560 4826
rect 56508 4762 56560 4768
rect 56888 3806 56916 64846
rect 56980 56166 57008 126647
rect 56968 56160 57020 56166
rect 56968 56102 57020 56108
rect 57072 4146 57100 143647
rect 57060 4140 57112 4146
rect 57060 4082 57112 4088
rect 56876 3800 56928 3806
rect 56876 3742 56928 3748
rect 55496 3596 55548 3602
rect 55496 3538 55548 3544
rect 56048 3596 56100 3602
rect 56048 3538 56100 3544
rect 56060 480 56088 3538
rect 57164 2922 57192 158607
rect 57256 3262 57284 234087
rect 57334 230752 57390 230761
rect 57334 230687 57390 230696
rect 57348 230518 57376 230687
rect 57336 230512 57388 230518
rect 57336 230454 57388 230460
rect 57336 230376 57388 230382
rect 57336 230318 57388 230324
rect 57244 3256 57296 3262
rect 57244 3198 57296 3204
rect 57242 3088 57298 3097
rect 57242 3023 57298 3032
rect 57152 2916 57204 2922
rect 57152 2858 57204 2864
rect 57256 480 57284 3023
rect 57348 2854 57376 230318
rect 57440 3670 57468 248367
rect 57428 3664 57480 3670
rect 57428 3606 57480 3612
rect 57532 3194 57560 329190
rect 57520 3188 57572 3194
rect 57520 3130 57572 3136
rect 57624 2990 57652 413607
rect 57716 208434 57744 630634
rect 57808 483721 57836 700674
rect 72988 700398 73016 703520
rect 59268 700392 59320 700398
rect 59268 700334 59320 700340
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 59082 533352 59138 533361
rect 59082 533287 59138 533296
rect 57794 483712 57850 483721
rect 57794 483647 57850 483656
rect 58990 472152 59046 472161
rect 58990 472087 59046 472096
rect 57794 449032 57850 449041
rect 57794 448967 57850 448976
rect 57808 208554 57836 448967
rect 58898 405512 58954 405521
rect 58898 405447 58954 405456
rect 58806 376272 58862 376281
rect 58806 376207 58862 376216
rect 57886 332752 57942 332761
rect 57886 332687 57942 332696
rect 57900 329254 57928 332687
rect 57888 329248 57940 329254
rect 57888 329190 57940 329196
rect 57978 321192 58034 321201
rect 57978 321127 58034 321136
rect 57886 294672 57942 294681
rect 57886 294607 57942 294616
rect 57900 294030 57928 294607
rect 57888 294024 57940 294030
rect 57888 293966 57940 293972
rect 57886 236872 57942 236881
rect 57886 236807 57942 236816
rect 57900 230382 57928 236807
rect 57888 230376 57940 230382
rect 57888 230318 57940 230324
rect 57886 228032 57942 228041
rect 57886 227967 57942 227976
rect 57900 227798 57928 227967
rect 57888 227792 57940 227798
rect 57888 227734 57940 227740
rect 57886 225312 57942 225321
rect 57886 225247 57942 225256
rect 57900 225010 57928 225247
rect 57888 225004 57940 225010
rect 57888 224946 57940 224952
rect 57886 222592 57942 222601
rect 57886 222527 57942 222536
rect 57900 222222 57928 222527
rect 57888 222216 57940 222222
rect 57888 222158 57940 222164
rect 57886 219192 57942 219201
rect 57886 219127 57942 219136
rect 57900 218074 57928 219127
rect 57888 218068 57940 218074
rect 57888 218010 57940 218016
rect 57886 211032 57942 211041
rect 57886 210967 57942 210976
rect 57900 209846 57928 210967
rect 57888 209840 57940 209846
rect 57888 209782 57940 209788
rect 57796 208548 57848 208554
rect 57796 208490 57848 208496
rect 57716 208406 57928 208434
rect 57704 208344 57756 208350
rect 57704 208286 57756 208292
rect 57796 208344 57848 208350
rect 57796 208286 57848 208292
rect 57716 207641 57744 208286
rect 57702 207632 57758 207641
rect 57702 207567 57758 207576
rect 57702 204912 57758 204921
rect 57702 204847 57758 204856
rect 57716 204338 57744 204847
rect 57704 204332 57756 204338
rect 57704 204274 57756 204280
rect 57702 196072 57758 196081
rect 57702 196007 57704 196016
rect 57756 196007 57758 196016
rect 57704 195978 57756 195984
rect 57704 194540 57756 194546
rect 57704 194482 57756 194488
rect 57716 193361 57744 194482
rect 57702 193352 57758 193361
rect 57702 193287 57758 193296
rect 57704 187672 57756 187678
rect 57704 187614 57756 187620
rect 57716 187241 57744 187614
rect 57702 187232 57758 187241
rect 57702 187167 57758 187176
rect 57702 184512 57758 184521
rect 57702 184447 57758 184456
rect 57716 183598 57744 184447
rect 57704 183592 57756 183598
rect 57704 183534 57756 183540
rect 57702 181792 57758 181801
rect 57702 181727 57758 181736
rect 57716 180878 57744 181727
rect 57704 180872 57756 180878
rect 57704 180814 57756 180820
rect 57702 172952 57758 172961
rect 57702 172887 57758 172896
rect 57716 172582 57744 172887
rect 57704 172576 57756 172582
rect 57704 172518 57756 172524
rect 57808 172514 57836 208286
rect 57900 202201 57928 208406
rect 57886 202192 57942 202201
rect 57886 202127 57942 202136
rect 57886 175672 57942 175681
rect 57886 175607 57942 175616
rect 57796 172508 57848 172514
rect 57796 172450 57848 172456
rect 57900 172394 57928 175607
rect 57716 172366 57928 172394
rect 57716 3058 57744 172366
rect 57796 172304 57848 172310
rect 57796 172246 57848 172252
rect 57808 3126 57836 172246
rect 57888 171080 57940 171086
rect 57888 171022 57940 171028
rect 57900 170241 57928 171022
rect 57886 170232 57942 170241
rect 57886 170167 57942 170176
rect 57886 166832 57942 166841
rect 57886 166767 57942 166776
rect 57900 165646 57928 166767
rect 57888 165640 57940 165646
rect 57888 165582 57940 165588
rect 57886 164112 57942 164121
rect 57886 164047 57942 164056
rect 57900 162926 57928 164047
rect 57888 162920 57940 162926
rect 57888 162862 57940 162868
rect 57888 155916 57940 155922
rect 57888 155858 57940 155864
rect 57900 155281 57928 155858
rect 57886 155272 57942 155281
rect 57886 155207 57942 155216
rect 57886 152552 57942 152561
rect 57886 152487 57942 152496
rect 57900 151842 57928 152487
rect 57888 151836 57940 151842
rect 57888 151778 57940 151784
rect 57886 149832 57942 149841
rect 57886 149767 57942 149776
rect 57900 149122 57928 149767
rect 57888 149116 57940 149122
rect 57888 149058 57940 149064
rect 57886 147112 57942 147121
rect 57886 147047 57942 147056
rect 57900 146334 57928 147047
rect 57888 146328 57940 146334
rect 57888 146270 57940 146276
rect 57886 140992 57942 141001
rect 57886 140927 57942 140936
rect 57900 140826 57928 140927
rect 57888 140820 57940 140826
rect 57888 140762 57940 140768
rect 57886 135552 57942 135561
rect 57886 135487 57942 135496
rect 57900 135318 57928 135487
rect 57888 135312 57940 135318
rect 57888 135254 57940 135260
rect 57886 132152 57942 132161
rect 57886 132087 57942 132096
rect 57900 131170 57928 132087
rect 57888 131164 57940 131170
rect 57888 131106 57940 131112
rect 57886 129432 57942 129441
rect 57886 129367 57942 129376
rect 57900 128382 57928 129367
rect 57888 128376 57940 128382
rect 57888 128318 57940 128324
rect 57886 123312 57942 123321
rect 57886 123247 57942 123256
rect 57900 122874 57928 123247
rect 57888 122868 57940 122874
rect 57888 122810 57940 122816
rect 57886 120592 57942 120601
rect 57886 120527 57942 120536
rect 57900 120154 57928 120527
rect 57888 120148 57940 120154
rect 57888 120090 57940 120096
rect 57886 117872 57942 117881
rect 57886 117807 57942 117816
rect 57900 117366 57928 117807
rect 57888 117360 57940 117366
rect 57888 117302 57940 117308
rect 57886 115152 57942 115161
rect 57886 115087 57942 115096
rect 57900 114578 57928 115087
rect 57888 114572 57940 114578
rect 57888 114514 57940 114520
rect 57888 107636 57940 107642
rect 57888 107578 57940 107584
rect 57900 106321 57928 107578
rect 57886 106312 57942 106321
rect 57886 106247 57942 106256
rect 57888 100700 57940 100706
rect 57888 100642 57940 100648
rect 57900 100201 57928 100642
rect 57886 100192 57942 100201
rect 57886 100127 57942 100136
rect 57886 94752 57942 94761
rect 57886 94687 57942 94696
rect 57900 93906 57928 94687
rect 57888 93900 57940 93906
rect 57888 93842 57940 93848
rect 57886 88632 57942 88641
rect 57886 88567 57942 88576
rect 57900 86018 57928 88567
rect 57888 86012 57940 86018
rect 57888 85954 57940 85960
rect 57886 85912 57942 85921
rect 57886 85847 57942 85856
rect 57900 85610 57928 85847
rect 57888 85604 57940 85610
rect 57888 85546 57940 85552
rect 57888 85468 57940 85474
rect 57888 85410 57940 85416
rect 57900 4078 57928 85410
rect 57992 16574 58020 321127
rect 58714 286512 58770 286521
rect 58714 286447 58770 286456
rect 58622 257272 58678 257281
rect 58622 257207 58678 257216
rect 58530 245712 58586 245721
rect 58530 245647 58586 245656
rect 58438 97472 58494 97481
rect 58438 97407 58494 97416
rect 58346 91352 58402 91361
rect 58346 91287 58402 91296
rect 58254 83192 58310 83201
rect 58254 83127 58310 83136
rect 58162 74352 58218 74361
rect 58162 74287 58218 74296
rect 58070 68232 58126 68241
rect 58070 68167 58126 68176
rect 58084 61810 58112 68167
rect 58072 61804 58124 61810
rect 58072 61746 58124 61752
rect 58176 56506 58204 74287
rect 58164 56500 58216 56506
rect 58164 56442 58216 56448
rect 58268 56370 58296 83127
rect 58256 56364 58308 56370
rect 58256 56306 58308 56312
rect 58360 28286 58388 91287
rect 58452 61538 58480 97407
rect 58440 61532 58492 61538
rect 58440 61474 58492 61480
rect 58544 60926 58572 245647
rect 58636 61334 58664 257207
rect 58624 61328 58676 61334
rect 58624 61270 58676 61276
rect 58532 60920 58584 60926
rect 58532 60862 58584 60868
rect 58348 28280 58400 28286
rect 58348 28222 58400 28228
rect 57992 16546 58480 16574
rect 57888 4072 57940 4078
rect 57888 4014 57940 4020
rect 57796 3120 57848 3126
rect 57796 3062 57848 3068
rect 57704 3052 57756 3058
rect 57704 2994 57756 3000
rect 57612 2984 57664 2990
rect 57612 2926 57664 2932
rect 57336 2848 57388 2854
rect 57336 2790 57388 2796
rect 58452 480 58480 16546
rect 58728 4486 58756 286447
rect 58820 5234 58848 376207
rect 58912 6186 58940 405447
rect 59004 61742 59032 472087
rect 58992 61736 59044 61742
rect 58992 61678 59044 61684
rect 59096 58682 59124 533287
rect 59174 501392 59230 501401
rect 59174 501327 59230 501336
rect 59084 58676 59136 58682
rect 59084 58618 59136 58624
rect 58900 6180 58952 6186
rect 58900 6122 58952 6128
rect 59188 5302 59216 501327
rect 59280 138281 59308 700334
rect 89180 697610 89208 703520
rect 92388 700800 92440 700806
rect 92388 700742 92440 700748
rect 89168 697604 89220 697610
rect 89168 697546 89220 697552
rect 89628 696992 89680 696998
rect 89628 696934 89680 696940
rect 89640 547874 89668 696934
rect 89456 547846 89668 547874
rect 80612 543312 80664 543318
rect 80612 543254 80664 543260
rect 61292 543176 61344 543182
rect 61292 543118 61344 543124
rect 78036 543176 78088 543182
rect 78036 543118 78088 543124
rect 61304 539852 61332 543118
rect 64512 543108 64564 543114
rect 64512 543050 64564 543056
rect 64524 539852 64552 543050
rect 67088 542496 67140 542502
rect 67088 542438 67140 542444
rect 67100 539852 67128 542438
rect 69664 542428 69716 542434
rect 69664 542370 69716 542376
rect 69676 539852 69704 542370
rect 78048 539852 78076 543118
rect 80624 539852 80652 543254
rect 89456 539866 89484 547846
rect 92400 543590 92428 700742
rect 91560 543584 91612 543590
rect 91560 543526 91612 543532
rect 92388 543584 92440 543590
rect 92388 543526 92440 543532
rect 89010 539838 89484 539866
rect 91572 539852 91600 543526
rect 94780 543244 94832 543250
rect 94780 543186 94832 543192
rect 94792 539852 94820 543186
rect 99932 543040 99984 543046
rect 99932 542982 99984 542988
rect 97356 542700 97408 542706
rect 97356 542642 97408 542648
rect 97368 539852 97396 542642
rect 99944 539852 99972 542982
rect 102508 542972 102560 542978
rect 102508 542914 102560 542920
rect 102520 539852 102548 542914
rect 104912 540326 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 122748 700664 122800 700670
rect 122748 700606 122800 700612
rect 122760 543590 122788 700606
rect 137848 700602 137876 703520
rect 144828 700868 144880 700874
rect 144828 700810 144880 700816
rect 137836 700596 137888 700602
rect 137836 700538 137888 700544
rect 136548 700392 136600 700398
rect 136548 700334 136600 700340
rect 136560 547874 136588 700334
rect 136376 547846 136588 547874
rect 121828 543584 121880 543590
rect 121828 543526 121880 543532
rect 122748 543584 122800 543590
rect 122748 543526 122800 543532
rect 132774 543552 132830 543561
rect 108304 543244 108356 543250
rect 108304 543186 108356 543192
rect 104900 540320 104952 540326
rect 104900 540262 104952 540268
rect 108316 539852 108344 543186
rect 113454 542600 113510 542609
rect 113454 542535 113510 542544
rect 113468 539852 113496 542535
rect 121840 539852 121868 543526
rect 132774 543487 132830 543496
rect 130200 542564 130252 542570
rect 130200 542506 130252 542512
rect 130212 539852 130240 542506
rect 132788 539852 132816 543487
rect 136376 539866 136404 547846
rect 144840 542570 144868 700810
rect 154132 700738 154160 703520
rect 170324 700874 170352 703520
rect 170312 700868 170364 700874
rect 170312 700810 170364 700816
rect 202800 700806 202828 703520
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 172428 700732 172480 700738
rect 172428 700674 172480 700680
rect 158628 616888 158680 616894
rect 158628 616830 158680 616836
rect 158640 543590 158668 616830
rect 164148 590708 164200 590714
rect 164148 590650 164200 590656
rect 164160 543590 164188 590650
rect 172440 543590 172468 700674
rect 218992 699825 219020 703520
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 218978 699816 219034 699825
rect 218978 699751 219034 699760
rect 267660 697678 267688 703520
rect 283852 700670 283880 703520
rect 300136 700738 300164 703520
rect 300124 700732 300176 700738
rect 300124 700674 300176 700680
rect 283840 700664 283892 700670
rect 283840 700606 283892 700612
rect 305000 700596 305052 700602
rect 305000 700538 305052 700544
rect 266360 697672 266412 697678
rect 266360 697614 266412 697620
rect 267648 697672 267700 697678
rect 267648 697614 267700 697620
rect 226798 543688 226854 543697
rect 226798 543623 226854 543632
rect 157892 543584 157944 543590
rect 157892 543526 157944 543532
rect 158628 543584 158680 543590
rect 158628 543526 158680 543532
rect 163044 543584 163096 543590
rect 163044 543526 163096 543532
rect 164148 543584 164200 543590
rect 164148 543526 164200 543532
rect 171416 543584 171468 543590
rect 171416 543526 171468 543532
rect 172428 543584 172480 543590
rect 172428 543526 172480 543532
rect 146942 542872 146998 542881
rect 146942 542807 146998 542816
rect 143724 542564 143776 542570
rect 143724 542506 143776 542512
rect 144828 542564 144880 542570
rect 144828 542506 144880 542512
rect 138570 542464 138626 542473
rect 138570 542399 138626 542408
rect 136022 539838 136404 539866
rect 138584 539852 138612 542399
rect 141424 539912 141476 539918
rect 141174 539860 141424 539866
rect 141174 539854 141476 539860
rect 141174 539838 141464 539854
rect 143736 539852 143764 542506
rect 146956 539852 146984 542807
rect 149518 542600 149574 542609
rect 149518 542535 149574 542544
rect 149532 539852 149560 542535
rect 152096 541000 152148 541006
rect 152096 540942 152148 540948
rect 152108 539852 152136 540942
rect 157904 539852 157932 543526
rect 163056 539852 163084 543526
rect 168838 543144 168894 543153
rect 168838 543079 168894 543088
rect 166262 543008 166318 543017
rect 166262 542943 166318 542952
rect 166276 539852 166304 542943
rect 168852 539852 168880 543079
rect 171428 539852 171456 543526
rect 179786 543416 179842 543425
rect 179786 543351 179842 543360
rect 173992 543312 174044 543318
rect 173992 543254 174044 543260
rect 174004 539852 174032 543254
rect 177210 542464 177266 542473
rect 177210 542399 177266 542408
rect 177224 539852 177252 542399
rect 179800 539852 179828 543351
rect 199108 542904 199160 542910
rect 199108 542846 199160 542852
rect 182364 542700 182416 542706
rect 182364 542642 182416 542648
rect 182376 539852 182404 542642
rect 190734 542464 190790 542473
rect 190734 542399 190790 542408
rect 185610 539850 185992 539866
rect 188186 539850 188568 539866
rect 190748 539852 190776 542399
rect 196532 541136 196584 541142
rect 196532 541078 196584 541084
rect 193680 539980 193732 539986
rect 193680 539922 193732 539928
rect 193692 539866 193720 539922
rect 185610 539844 186004 539850
rect 185610 539838 185952 539844
rect 188186 539844 188580 539850
rect 188186 539838 188528 539844
rect 185952 539786 186004 539792
rect 193338 539838 193720 539866
rect 196544 539852 196572 541078
rect 199120 539852 199148 542846
rect 204260 542836 204312 542842
rect 204260 542778 204312 542784
rect 201960 539980 202012 539986
rect 201960 539922 202012 539928
rect 201972 539866 202000 539922
rect 201710 539838 202000 539866
rect 204272 539852 204300 542778
rect 210054 542600 210110 542609
rect 210054 542535 210110 542544
rect 207204 539980 207256 539986
rect 207204 539922 207256 539928
rect 207216 539866 207244 539922
rect 207216 539838 207506 539866
rect 210068 539852 210096 542535
rect 215206 541240 215262 541249
rect 215206 541175 215262 541184
rect 212632 541068 212684 541074
rect 212632 541010 212684 541016
rect 212644 539852 212672 541010
rect 215220 539852 215248 541175
rect 218704 539980 218756 539986
rect 218704 539922 218756 539928
rect 218716 539866 218744 539922
rect 218454 539838 218744 539866
rect 226812 539852 226840 543623
rect 259644 542904 259696 542910
rect 259644 542846 259696 542852
rect 248696 542836 248748 542842
rect 248696 542778 248748 542784
rect 231950 542464 232006 542473
rect 231950 542399 232006 542408
rect 229744 539980 229796 539986
rect 229744 539922 229796 539928
rect 229756 539866 229784 539922
rect 229402 539838 229784 539866
rect 231964 539852 231992 542399
rect 237748 541272 237800 541278
rect 237748 541214 237800 541220
rect 234436 539980 234488 539986
rect 234436 539922 234488 539928
rect 234448 539866 234476 539922
rect 234448 539838 234554 539866
rect 237760 539852 237788 541214
rect 245384 540048 245436 540054
rect 245384 539990 245436 539996
rect 245396 539866 245424 539990
rect 245396 539838 245502 539866
rect 248708 539852 248736 542778
rect 251270 542600 251326 542609
rect 251270 542535 251326 542544
rect 251284 539852 251312 542535
rect 257066 542464 257122 542473
rect 257066 542399 257122 542408
rect 257080 539852 257108 542399
rect 259656 539852 259684 542846
rect 266372 541686 266400 697614
rect 281540 579692 281592 579698
rect 281540 579634 281592 579640
rect 275744 542768 275796 542774
rect 275744 542710 275796 542716
rect 266360 541680 266412 541686
rect 266360 541622 266412 541628
rect 264796 541204 264848 541210
rect 264796 541146 264848 541152
rect 262220 540116 262272 540122
rect 262220 540058 262272 540064
rect 262232 539852 262260 540058
rect 264808 539852 264836 541146
rect 268384 540048 268436 540054
rect 268384 539990 268436 539996
rect 272892 540048 272944 540054
rect 272892 539990 272944 539996
rect 268396 539866 268424 539990
rect 268042 539838 268424 539866
rect 272904 539866 272932 539990
rect 272904 539838 273194 539866
rect 275756 539852 275784 542710
rect 281552 539852 281580 579634
rect 305012 557534 305040 700538
rect 332520 700534 332548 703520
rect 348804 700534 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 305012 557506 305592 557534
rect 292486 543280 292542 543289
rect 292486 543215 292542 543224
rect 287152 540048 287204 540054
rect 287152 539990 287204 539996
rect 289820 540048 289872 540054
rect 289820 539990 289872 539996
rect 287164 539866 287192 539990
rect 289832 539866 289860 539990
rect 287164 539838 287362 539866
rect 289832 539838 289938 539866
rect 292500 539852 292528 543215
rect 300860 540116 300912 540122
rect 300860 540058 300912 540064
rect 303436 540116 303488 540122
rect 303436 540058 303488 540064
rect 295248 540048 295300 540054
rect 295248 539990 295300 539996
rect 295260 539866 295288 539990
rect 295090 539838 295288 539866
rect 300872 539852 300900 540058
rect 303448 539852 303476 540058
rect 305564 539866 305592 557506
rect 347226 543144 347282 543153
rect 347226 543079 347282 543088
rect 311806 543008 311862 543017
rect 311806 542943 311862 542952
rect 305564 539838 306038 539866
rect 311820 539852 311848 542943
rect 325332 542768 325384 542774
rect 325332 542710 325384 542716
rect 336278 542736 336334 542745
rect 320180 540116 320232 540122
rect 320180 540058 320232 540064
rect 322756 540116 322808 540122
rect 322756 540058 322808 540064
rect 320192 539852 320220 540058
rect 322768 539852 322796 540058
rect 325344 539852 325372 542710
rect 336278 542671 336334 542680
rect 333704 542632 333756 542638
rect 333704 542574 333756 542580
rect 328552 540116 328604 540122
rect 328552 540058 328604 540064
rect 328564 539852 328592 540058
rect 333716 539852 333744 542574
rect 336292 539852 336320 542671
rect 344652 541408 344704 541414
rect 344652 541350 344704 541356
rect 339500 540116 339552 540122
rect 339500 540058 339552 540064
rect 339512 539852 339540 540058
rect 344664 539852 344692 541350
rect 347240 539852 347268 543079
rect 358818 542872 358874 542881
rect 358818 542807 358874 542816
rect 353022 542600 353078 542609
rect 353022 542535 353078 542544
rect 353036 539852 353064 542535
rect 355600 540116 355652 540122
rect 355600 540058 355652 540064
rect 355612 539852 355640 540058
rect 358832 539852 358860 542807
rect 364352 540258 364380 702406
rect 397472 700466 397500 703520
rect 413664 700466 413692 703520
rect 429856 700602 429884 703520
rect 439504 700664 439556 700670
rect 439504 700606 439556 700612
rect 429844 700596 429896 700602
rect 429844 700538 429896 700544
rect 397460 700460 397512 700466
rect 397460 700402 397512 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 439412 670744 439464 670750
rect 439412 670686 439464 670692
rect 427084 543380 427136 543386
rect 427084 543322 427136 543328
rect 418712 543108 418764 543114
rect 418712 543050 418764 543056
rect 407764 543040 407816 543046
rect 407764 542982 407816 542988
rect 410982 543008 411038 543017
rect 369768 542972 369820 542978
rect 369768 542914 369820 542920
rect 366546 542600 366602 542609
rect 366546 542535 366602 542544
rect 364340 540252 364392 540258
rect 364340 540194 364392 540200
rect 363972 540116 364024 540122
rect 363972 540058 364024 540064
rect 363984 539852 364012 540058
rect 366560 539852 366588 542535
rect 369780 539852 369808 542914
rect 391662 542872 391718 542881
rect 391662 542807 391718 542816
rect 380714 542736 380770 542745
rect 380714 542671 380770 542680
rect 374920 541612 374972 541618
rect 374920 541554 374972 541560
rect 372344 541544 372396 541550
rect 372344 541486 372396 541492
rect 372356 539852 372384 541486
rect 374932 539852 374960 541554
rect 380728 539852 380756 542671
rect 391676 539852 391704 542807
rect 405188 542632 405240 542638
rect 396814 542600 396870 542609
rect 405188 542574 405240 542580
rect 396814 542535 396870 542544
rect 396828 539852 396856 542535
rect 400036 541476 400088 541482
rect 400036 541418 400088 541424
rect 400048 539852 400076 541418
rect 405200 539852 405228 542574
rect 407776 539852 407804 542982
rect 410982 542943 411038 542952
rect 410996 539852 411024 542943
rect 413560 540184 413612 540190
rect 413560 540126 413612 540132
rect 416136 540184 416188 540190
rect 416136 540126 416188 540132
rect 413572 539852 413600 540126
rect 416148 539852 416176 540126
rect 418724 539852 418752 543050
rect 421932 541340 421984 541346
rect 421932 541282 421984 541288
rect 421944 539852 421972 541282
rect 424508 540184 424560 540190
rect 424508 540126 424560 540132
rect 424520 539852 424548 540126
rect 427096 539852 427124 543322
rect 430304 542496 430356 542502
rect 430304 542438 430356 542444
rect 430316 539852 430344 542438
rect 432880 542428 432932 542434
rect 432880 542370 432932 542376
rect 432892 539852 432920 542370
rect 188528 539786 188580 539792
rect 110906 539714 111288 539730
rect 110906 539708 111300 539714
rect 110906 539702 111248 539708
rect 111248 539650 111300 539656
rect 86776 539640 86828 539646
rect 72606 539608 72662 539617
rect 72266 539566 72606 539594
rect 75642 539608 75698 539617
rect 75486 539566 75642 539594
rect 72606 539543 72662 539552
rect 83858 539578 84056 539594
rect 86434 539588 86776 539594
rect 106094 539608 106150 539617
rect 86434 539582 86828 539588
rect 83858 539572 84068 539578
rect 83858 539566 84016 539572
rect 75642 539543 75698 539552
rect 86434 539566 86816 539582
rect 105754 539566 106094 539594
rect 106094 539543 106150 539552
rect 116306 539608 116362 539617
rect 119526 539608 119582 539617
rect 116362 539566 116702 539594
rect 119278 539566 119526 539594
rect 116306 539543 116362 539552
rect 125322 539608 125378 539617
rect 125074 539566 125322 539594
rect 119526 539543 119582 539552
rect 125322 539543 125378 539552
rect 127346 539608 127402 539617
rect 155590 539608 155646 539617
rect 127402 539566 127650 539594
rect 155342 539566 155590 539594
rect 127346 539543 127402 539552
rect 220634 539608 220690 539617
rect 160494 539578 160784 539594
rect 160494 539572 160796 539578
rect 160494 539566 160744 539572
rect 155590 539543 155646 539552
rect 84016 539514 84068 539520
rect 243174 539608 243230 539617
rect 220690 539566 221030 539594
rect 242926 539566 243174 539594
rect 220634 539543 220690 539552
rect 243174 539543 243230 539552
rect 253570 539608 253626 539617
rect 283838 539608 283894 539617
rect 253626 539566 253874 539594
rect 253570 539543 253626 539552
rect 314106 539608 314162 539617
rect 283894 539566 284142 539594
rect 283838 539543 283894 539552
rect 330850 539608 330906 539617
rect 314162 539566 314410 539594
rect 314106 539543 314162 539552
rect 341706 539608 341762 539617
rect 330906 539566 331154 539594
rect 330850 539543 330906 539552
rect 361026 539608 361082 539617
rect 341762 539566 342102 539594
rect 341706 539543 341762 539552
rect 377310 539608 377366 539617
rect 361082 539566 361422 539594
rect 361026 539543 361082 539552
rect 382922 539608 382978 539617
rect 377366 539566 377522 539594
rect 377310 539543 377366 539552
rect 385498 539608 385554 539617
rect 382978 539566 383318 539594
rect 382922 539543 382978 539552
rect 388810 539608 388866 539617
rect 385554 539566 385894 539594
rect 385498 539543 385554 539552
rect 393962 539608 394018 539617
rect 388866 539566 389114 539594
rect 388810 539543 388866 539552
rect 402242 539608 402298 539617
rect 394018 539566 394266 539594
rect 393962 539543 394018 539552
rect 402298 539566 402638 539594
rect 438058 539578 438440 539594
rect 438058 539572 438452 539578
rect 438058 539566 438400 539572
rect 402242 539543 402298 539552
rect 160744 539514 160796 539520
rect 438400 539514 438452 539520
rect 435180 539504 435232 539510
rect 60646 539472 60702 539481
rect 60646 539407 60648 539416
rect 60700 539407 60702 539416
rect 223486 539472 223542 539481
rect 240230 539472 240286 539481
rect 223542 539430 223606 539458
rect 223486 539407 223542 539416
rect 270314 539472 270370 539481
rect 240286 539430 240350 539458
rect 240230 539407 240286 539416
rect 278870 539472 278926 539481
rect 270370 539430 270618 539458
rect 270314 539407 270370 539416
rect 298190 539472 298246 539481
rect 278926 539430 278990 539458
rect 278870 539407 278926 539416
rect 309138 539472 309194 539481
rect 298246 539430 298310 539458
rect 298190 539407 298246 539416
rect 350354 539472 350410 539481
rect 309194 539430 309258 539458
rect 309138 539407 309194 539416
rect 350410 539430 350474 539458
rect 435232 539452 435482 539458
rect 435180 539446 435482 539452
rect 435192 539430 435482 539446
rect 350354 539407 350410 539416
rect 60648 539378 60700 539384
rect 316972 539238 317000 539308
rect 316960 539232 317012 539238
rect 316960 539174 317012 539180
rect 59820 537940 59872 537946
rect 59820 537882 59872 537888
rect 59832 536625 59860 537882
rect 59818 536616 59874 536625
rect 59818 536551 59874 536560
rect 59358 497992 59414 498001
rect 59358 497927 59414 497936
rect 59266 138272 59322 138281
rect 59266 138207 59322 138216
rect 59266 109032 59322 109041
rect 59266 108967 59322 108976
rect 59280 60382 59308 108967
rect 59268 60376 59320 60382
rect 59268 60318 59320 60324
rect 59372 5370 59400 497927
rect 59450 425912 59506 425921
rect 59450 425847 59506 425856
rect 59360 5364 59412 5370
rect 59360 5306 59412 5312
rect 59176 5296 59228 5302
rect 59176 5238 59228 5244
rect 58808 5228 58860 5234
rect 58808 5170 58860 5176
rect 59464 4690 59492 425847
rect 59542 318472 59598 318481
rect 59542 318407 59598 318416
rect 59556 5846 59584 318407
rect 59634 306232 59690 306241
rect 59634 306167 59690 306176
rect 59648 54806 59676 306167
rect 439424 152402 439452 670686
rect 439516 445913 439544 700606
rect 440424 700596 440476 700602
rect 440424 700538 440476 700544
rect 439872 700528 439924 700534
rect 439872 700470 439924 700476
rect 439780 700460 439832 700466
rect 439780 700402 439832 700408
rect 439596 543244 439648 543250
rect 439596 543186 439648 543192
rect 439502 445904 439558 445913
rect 439502 445839 439558 445848
rect 439502 438968 439558 438977
rect 439502 438903 439558 438912
rect 439516 152522 439544 438903
rect 439608 152522 439636 543186
rect 439688 542428 439740 542434
rect 439688 542370 439740 542376
rect 439700 171134 439728 542370
rect 439792 387705 439820 700402
rect 439884 495145 439912 700470
rect 440332 656940 440384 656946
rect 440332 656882 440384 656888
rect 440240 539504 440292 539510
rect 440240 539446 440292 539452
rect 439962 537976 440018 537985
rect 439962 537911 440018 537920
rect 439976 537878 440004 537911
rect 439964 537872 440016 537878
rect 439964 537814 440016 537820
rect 439870 495136 439926 495145
rect 439870 495071 439926 495080
rect 439778 387696 439834 387705
rect 439778 387631 439834 387640
rect 439700 171106 439912 171134
rect 439504 152516 439556 152522
rect 439504 152458 439556 152464
rect 439596 152516 439648 152522
rect 439596 152458 439648 152464
rect 439502 152416 439558 152425
rect 439424 152374 439502 152402
rect 439502 152351 439558 152360
rect 439504 152312 439556 152318
rect 439504 152254 439556 152260
rect 439596 152312 439648 152318
rect 439596 152254 439648 152260
rect 59726 111752 59782 111761
rect 59726 111687 59782 111696
rect 59740 58546 59768 111687
rect 59818 79792 59874 79801
rect 59818 79727 59874 79736
rect 59832 74534 59860 79727
rect 59832 74506 59952 74534
rect 59818 62792 59874 62801
rect 59818 62727 59874 62736
rect 59728 58540 59780 58546
rect 59728 58482 59780 58488
rect 59832 56302 59860 62727
rect 59924 60450 59952 74506
rect 439516 73234 439544 152254
rect 439504 73228 439556 73234
rect 439504 73170 439556 73176
rect 439502 73128 439558 73137
rect 439424 73086 439502 73114
rect 176660 60648 176712 60654
rect 176660 60590 176712 60596
rect 200028 60648 200080 60654
rect 200028 60590 200080 60596
rect 160100 60580 160152 60586
rect 160100 60522 160152 60528
rect 168288 60580 168340 60586
rect 168288 60522 168340 60528
rect 59912 60444 59964 60450
rect 59912 60386 59964 60392
rect 135260 60444 135312 60450
rect 135260 60386 135312 60392
rect 143540 60444 143592 60450
rect 143540 60386 143592 60392
rect 149152 60444 149204 60450
rect 149152 60386 149204 60392
rect 151728 60444 151780 60450
rect 151728 60386 151780 60392
rect 67640 60376 67692 60382
rect 67640 60318 67692 60324
rect 80060 60376 80112 60382
rect 80060 60318 80112 60324
rect 122748 60376 122800 60382
rect 122748 60318 122800 60324
rect 60016 57798 60044 60044
rect 60004 57792 60056 57798
rect 60004 57734 60056 57740
rect 62592 57730 62620 60044
rect 62580 57724 62632 57730
rect 62580 57666 62632 57672
rect 63316 57724 63368 57730
rect 63316 57666 63368 57672
rect 59820 56296 59872 56302
rect 59820 56238 59872 56244
rect 59636 54800 59688 54806
rect 59636 54742 59688 54748
rect 62028 50448 62080 50454
rect 62028 50390 62080 50396
rect 59544 5840 59596 5846
rect 59544 5782 59596 5788
rect 59452 4684 59504 4690
rect 59452 4626 59504 4632
rect 58716 4480 58768 4486
rect 58716 4422 58768 4428
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 59648 480 59676 3538
rect 60830 2816 60886 2825
rect 60830 2751 60886 2760
rect 60844 480 60872 2751
rect 62040 480 62068 50390
rect 63328 5098 63356 57666
rect 63408 57180 63460 57186
rect 63408 57122 63460 57128
rect 63316 5092 63368 5098
rect 63316 5034 63368 5040
rect 63420 3482 63448 57122
rect 65168 56710 65196 60044
rect 65156 56704 65208 56710
rect 65156 56646 65208 56652
rect 66076 56704 66128 56710
rect 66076 56646 66128 56652
rect 66088 5030 66116 56646
rect 66168 56228 66220 56234
rect 66168 56170 66220 56176
rect 66076 5024 66128 5030
rect 66076 4966 66128 4972
rect 66180 3942 66208 56170
rect 67652 16574 67680 60318
rect 67744 57730 67772 60044
rect 70412 60030 70978 60058
rect 69756 57792 69808 57798
rect 69756 57734 69808 57740
rect 67732 57724 67784 57730
rect 67732 57666 67784 57672
rect 68928 57724 68980 57730
rect 68928 57666 68980 57672
rect 67652 16546 67956 16574
rect 65524 3936 65576 3942
rect 64326 3904 64382 3913
rect 65524 3878 65576 3884
rect 66168 3936 66220 3942
rect 66168 3878 66220 3884
rect 64326 3839 64382 3848
rect 63236 3454 63448 3482
rect 63236 480 63264 3454
rect 64340 480 64368 3839
rect 65536 480 65564 3878
rect 66718 2816 66774 2825
rect 66718 2751 66774 2760
rect 66732 480 66760 2751
rect 67928 480 67956 16546
rect 68940 4758 68968 57666
rect 69768 45554 69796 57734
rect 69676 45526 69796 45554
rect 69112 6860 69164 6866
rect 69112 6802 69164 6808
rect 68928 4752 68980 4758
rect 68928 4694 68980 4700
rect 69124 480 69152 6802
rect 69676 6254 69704 45526
rect 69664 6248 69716 6254
rect 69664 6190 69716 6196
rect 70308 4004 70360 4010
rect 70308 3946 70360 3952
rect 70320 480 70348 3946
rect 70412 3942 70440 60030
rect 73540 57866 73568 60044
rect 73528 57860 73580 57866
rect 73528 57802 73580 57808
rect 74448 57860 74500 57866
rect 74448 57802 74500 57808
rect 74460 6254 74488 57802
rect 76116 56914 76144 60044
rect 77208 58812 77260 58818
rect 77208 58754 77260 58760
rect 76104 56908 76156 56914
rect 76104 56850 76156 56856
rect 74448 6248 74500 6254
rect 74448 6190 74500 6196
rect 77220 4146 77248 58754
rect 71504 4140 71556 4146
rect 71504 4082 71556 4088
rect 71688 4140 71740 4146
rect 71688 4082 71740 4088
rect 76196 4140 76248 4146
rect 76196 4082 76248 4088
rect 77208 4140 77260 4146
rect 77208 4082 77260 4088
rect 70400 3936 70452 3942
rect 70400 3878 70452 3884
rect 71516 480 71544 4082
rect 71596 3936 71648 3942
rect 71596 3878 71648 3884
rect 71608 2825 71636 3878
rect 71700 3097 71728 4082
rect 72608 4072 72660 4078
rect 72608 4014 72660 4020
rect 71686 3088 71742 3097
rect 71686 3023 71742 3032
rect 71594 2816 71650 2825
rect 71594 2751 71650 2760
rect 72620 480 72648 4014
rect 73802 3224 73858 3233
rect 73802 3159 73858 3168
rect 73816 480 73844 3159
rect 75000 2916 75052 2922
rect 75000 2858 75052 2864
rect 75012 480 75040 2858
rect 76208 480 76236 4082
rect 78588 3936 78640 3942
rect 78588 3878 78640 3884
rect 77392 2916 77444 2922
rect 77392 2858 77444 2864
rect 77404 480 77432 2858
rect 78600 480 78628 3878
rect 78692 3602 78720 60044
rect 79968 49020 80020 49026
rect 79968 48962 80020 48968
rect 78680 3596 78732 3602
rect 78680 3538 78732 3544
rect 79980 2774 80008 48962
rect 80072 16574 80100 60318
rect 82820 60308 82872 60314
rect 82820 60250 82872 60256
rect 99288 60308 99340 60314
rect 99288 60250 99340 60256
rect 81532 57724 81584 57730
rect 81532 57666 81584 57672
rect 81544 16574 81572 57666
rect 81912 57390 81940 60044
rect 81900 57384 81952 57390
rect 81900 57326 81952 57332
rect 80072 16546 80928 16574
rect 81544 16546 82124 16574
rect 79704 2746 80008 2774
rect 79704 480 79732 2746
rect 80900 480 80928 16546
rect 82096 480 82124 16546
rect 82832 3602 82860 60250
rect 84488 59362 84516 60044
rect 84476 59356 84528 59362
rect 84476 59298 84528 59304
rect 87064 57730 87092 60044
rect 87052 57724 87104 57730
rect 87052 57666 87104 57672
rect 89640 57390 89668 60044
rect 92860 57866 92888 60044
rect 92848 57860 92900 57866
rect 92848 57802 92900 57808
rect 89628 57384 89680 57390
rect 89628 57326 89680 57332
rect 95436 57322 95464 60044
rect 95424 57316 95476 57322
rect 95424 57258 95476 57264
rect 83464 56908 83516 56914
rect 83464 56850 83516 56856
rect 83476 13258 83504 56850
rect 98012 56778 98040 60044
rect 98000 56772 98052 56778
rect 98000 56714 98052 56720
rect 99196 56772 99248 56778
rect 99196 56714 99248 56720
rect 95148 50516 95200 50522
rect 95148 50458 95200 50464
rect 83464 13252 83516 13258
rect 83464 13194 83516 13200
rect 90364 6656 90416 6662
rect 90364 6598 90416 6604
rect 86868 6044 86920 6050
rect 86868 5986 86920 5992
rect 82820 3596 82872 3602
rect 82820 3538 82872 3544
rect 83280 3596 83332 3602
rect 83280 3538 83332 3544
rect 84476 3596 84528 3602
rect 84476 3538 84528 3544
rect 83292 480 83320 3538
rect 84488 480 84516 3538
rect 85672 2848 85724 2854
rect 85672 2790 85724 2796
rect 85684 480 85712 2790
rect 86880 480 86908 5986
rect 89168 2984 89220 2990
rect 89168 2926 89220 2932
rect 87972 2848 88024 2854
rect 87972 2790 88024 2796
rect 87984 480 88012 2790
rect 89180 480 89208 2926
rect 90376 480 90404 6598
rect 95160 3670 95188 50458
rect 99208 46918 99236 56714
rect 99196 46912 99248 46918
rect 99196 46854 99248 46860
rect 99300 3670 99328 60250
rect 101232 57798 101260 60044
rect 102232 57860 102284 57866
rect 102232 57802 102284 57808
rect 101220 57792 101272 57798
rect 101220 57734 101272 57740
rect 100668 57044 100720 57050
rect 100668 56986 100720 56992
rect 100680 3670 100708 56986
rect 102244 16574 102272 57802
rect 103808 57118 103836 60044
rect 106384 57798 106412 60044
rect 108960 59430 108988 60044
rect 108948 59424 109000 59430
rect 108948 59366 109000 59372
rect 112180 57798 112208 60044
rect 114756 59294 114784 60044
rect 114744 59288 114796 59294
rect 114744 59230 114796 59236
rect 104808 57792 104860 57798
rect 104808 57734 104860 57740
rect 106372 57792 106424 57798
rect 106372 57734 106424 57740
rect 112168 57792 112220 57798
rect 112168 57734 112220 57740
rect 112996 57792 113048 57798
rect 112996 57734 113048 57740
rect 103796 57112 103848 57118
rect 103796 57054 103848 57060
rect 102244 16546 103376 16574
rect 101036 5976 101088 5982
rect 101036 5918 101088 5924
rect 91560 3664 91612 3670
rect 91560 3606 91612 3612
rect 93952 3664 94004 3670
rect 93952 3606 94004 3612
rect 95148 3664 95200 3670
rect 95148 3606 95200 3612
rect 98644 3664 98696 3670
rect 98644 3606 98696 3612
rect 99288 3664 99340 3670
rect 99288 3606 99340 3612
rect 99840 3664 99892 3670
rect 99840 3606 99892 3612
rect 100668 3664 100720 3670
rect 100668 3606 100720 3612
rect 91572 480 91600 3606
rect 92754 2816 92810 2825
rect 92754 2751 92810 2760
rect 92768 480 92796 2751
rect 93964 480 93992 3606
rect 97448 3120 97500 3126
rect 97448 3062 97500 3068
rect 96252 3052 96304 3058
rect 96252 2994 96304 3000
rect 95148 2984 95200 2990
rect 95148 2926 95200 2932
rect 95160 480 95188 2926
rect 96264 480 96292 2994
rect 97460 480 97488 3062
rect 98656 480 98684 3606
rect 99852 480 99880 3606
rect 101048 480 101076 5918
rect 102232 3800 102284 3806
rect 102232 3742 102284 3748
rect 102244 480 102272 3742
rect 103348 480 103376 16546
rect 104820 6914 104848 57734
rect 111708 50584 111760 50590
rect 111708 50526 111760 50532
rect 111720 6914 111748 50526
rect 104544 6886 104848 6914
rect 111628 6886 111748 6914
rect 104544 480 104572 6886
rect 109314 4040 109370 4049
rect 109314 3975 109370 3984
rect 108118 3088 108174 3097
rect 105728 3052 105780 3058
rect 108118 3023 108174 3032
rect 105728 2994 105780 3000
rect 105740 480 105768 2994
rect 106922 2952 106978 2961
rect 106922 2887 106978 2896
rect 106936 480 106964 2887
rect 108132 480 108160 3023
rect 109328 480 109356 3975
rect 110510 2952 110566 2961
rect 110510 2887 110566 2896
rect 110524 480 110552 2887
rect 111628 480 111656 6886
rect 113008 5506 113036 57734
rect 113088 56908 113140 56914
rect 113088 56850 113140 56856
rect 112996 5500 113048 5506
rect 112996 5442 113048 5448
rect 113100 3482 113128 56850
rect 117332 56642 117360 60044
rect 119908 57322 119936 60044
rect 119896 57316 119948 57322
rect 119896 57258 119948 57264
rect 117320 56636 117372 56642
rect 117320 56578 117372 56584
rect 116400 6724 116452 6730
rect 116400 6666 116452 6672
rect 114008 5908 114060 5914
rect 114008 5850 114060 5856
rect 112824 3454 113128 3482
rect 112824 480 112852 3454
rect 114020 480 114048 5850
rect 115204 2984 115256 2990
rect 115204 2926 115256 2932
rect 115216 480 115244 2926
rect 116412 480 116440 6666
rect 117594 4040 117650 4049
rect 117594 3975 117650 3984
rect 117608 480 117636 3975
rect 122760 3806 122788 60318
rect 123128 57866 123156 60044
rect 123116 57860 123168 57866
rect 123116 57802 123168 57808
rect 125704 56982 125732 60044
rect 127912 60030 128294 60058
rect 127164 59900 127216 59906
rect 127164 59842 127216 59848
rect 125692 56976 125744 56982
rect 125692 56918 125744 56924
rect 126888 56976 126940 56982
rect 126888 56918 126940 56924
rect 123484 56636 123536 56642
rect 123484 56578 123536 56584
rect 123496 15910 123524 56578
rect 123484 15904 123536 15910
rect 123484 15846 123536 15852
rect 126796 11824 126848 11830
rect 126796 11766 126848 11772
rect 125508 10736 125560 10742
rect 125508 10678 125560 10684
rect 122288 3800 122340 3806
rect 122288 3742 122340 3748
rect 122748 3800 122800 3806
rect 122748 3742 122800 3748
rect 121092 3188 121144 3194
rect 121092 3130 121144 3136
rect 119896 3120 119948 3126
rect 118790 3088 118846 3097
rect 119896 3062 119948 3068
rect 118790 3023 118846 3032
rect 118804 480 118832 3023
rect 119908 480 119936 3062
rect 121104 480 121132 3130
rect 122300 480 122328 3742
rect 125520 3262 125548 10678
rect 126808 3262 126836 11766
rect 126900 7954 126928 56918
rect 126888 7948 126940 7954
rect 126888 7890 126940 7896
rect 127176 6914 127204 59842
rect 127912 57594 127940 60030
rect 131500 57798 131528 60044
rect 131488 57792 131540 57798
rect 131488 57734 131540 57740
rect 127900 57588 127952 57594
rect 127900 57530 127952 57536
rect 128268 57588 128320 57594
rect 128268 57530 128320 57536
rect 128280 6914 128308 57530
rect 134076 56982 134104 60044
rect 134064 56976 134116 56982
rect 134064 56918 134116 56924
rect 129648 56772 129700 56778
rect 129648 56714 129700 56720
rect 129660 6914 129688 56714
rect 135168 54732 135220 54738
rect 135168 54674 135220 54680
rect 132408 51944 132460 51950
rect 132408 51886 132460 51892
rect 129740 47592 129792 47598
rect 129740 47534 129792 47540
rect 129752 16574 129780 47534
rect 129752 16546 130608 16574
rect 126992 6886 127204 6914
rect 128188 6886 128308 6914
rect 129384 6886 129688 6914
rect 123484 3256 123536 3262
rect 123484 3198 123536 3204
rect 124680 3256 124732 3262
rect 124680 3198 124732 3204
rect 125508 3256 125560 3262
rect 125508 3198 125560 3204
rect 125876 3256 125928 3262
rect 125876 3198 125928 3204
rect 126796 3256 126848 3262
rect 126796 3198 126848 3204
rect 123496 480 123524 3198
rect 124692 480 124720 3198
rect 125888 480 125916 3198
rect 126992 480 127020 6886
rect 128188 480 128216 6886
rect 129384 480 129412 6886
rect 130580 480 130608 16546
rect 132420 3262 132448 51886
rect 132960 5160 133012 5166
rect 132960 5102 133012 5108
rect 131764 3256 131816 3262
rect 131764 3198 131816 3204
rect 132408 3256 132460 3262
rect 132408 3198 132460 3204
rect 131776 480 131804 3198
rect 132972 480 133000 5102
rect 135180 3262 135208 54674
rect 134156 3256 134208 3262
rect 134156 3198 134208 3204
rect 135168 3256 135220 3262
rect 135168 3198 135220 3204
rect 134168 480 134196 3198
rect 135272 480 135300 60386
rect 136652 57798 136680 60044
rect 136640 57792 136692 57798
rect 136640 57734 136692 57740
rect 139228 57662 139256 60044
rect 142448 57798 142476 60044
rect 142436 57792 142488 57798
rect 142436 57734 142488 57740
rect 143448 57792 143500 57798
rect 143448 57734 143500 57740
rect 139216 57656 139268 57662
rect 139216 57598 139268 57604
rect 140044 57656 140096 57662
rect 140044 57598 140096 57604
rect 140056 25566 140084 57598
rect 140044 25560 140096 25566
rect 140044 25502 140096 25508
rect 137926 21312 137982 21321
rect 137926 21247 137982 21256
rect 137940 6914 137968 21247
rect 139306 13016 139362 13025
rect 139306 12951 139362 12960
rect 137664 6886 137968 6914
rect 136456 4480 136508 4486
rect 136456 4422 136508 4428
rect 136468 480 136496 4422
rect 137664 480 137692 6886
rect 139320 3262 139348 12951
rect 142436 4616 142488 4622
rect 142436 4558 142488 4564
rect 141240 4548 141292 4554
rect 141240 4490 141292 4496
rect 140044 4480 140096 4486
rect 140044 4422 140096 4428
rect 138848 3256 138900 3262
rect 138848 3198 138900 3204
rect 139308 3256 139360 3262
rect 139308 3198 139360 3204
rect 138860 480 138888 3198
rect 140056 480 140084 4422
rect 141252 480 141280 4490
rect 142448 480 142476 4558
rect 143460 4554 143488 57734
rect 143448 4548 143500 4554
rect 143448 4490 143500 4496
rect 143552 480 143580 60386
rect 145024 57798 145052 60044
rect 145012 57792 145064 57798
rect 145012 57734 145064 57740
rect 146208 57792 146260 57798
rect 146208 57734 146260 57740
rect 144826 24168 144882 24177
rect 144826 24103 144882 24112
rect 144840 6914 144868 24103
rect 145930 11656 145986 11665
rect 145930 11591 145986 11600
rect 144748 6886 144868 6914
rect 144748 480 144776 6886
rect 145944 480 145972 11591
rect 146220 4622 146248 57734
rect 147128 8220 147180 8226
rect 147128 8162 147180 8168
rect 146208 4616 146260 4622
rect 146208 4558 146260 4564
rect 147140 480 147168 8162
rect 147600 7410 147628 60044
rect 148968 57792 149020 57798
rect 148968 57734 149020 57740
rect 147588 7404 147640 7410
rect 147588 7346 147640 7352
rect 148980 3330 149008 57734
rect 149164 16574 149192 60386
rect 150176 57050 150204 60044
rect 150164 57044 150216 57050
rect 150164 56986 150216 56992
rect 149164 16546 149560 16574
rect 148324 3324 148376 3330
rect 148324 3266 148376 3272
rect 148968 3324 149020 3330
rect 148968 3266 149020 3272
rect 148336 480 148364 3266
rect 149532 480 149560 16546
rect 151740 3330 151768 60386
rect 153212 60030 153410 60058
rect 153016 5840 153068 5846
rect 153016 5782 153068 5788
rect 151820 5432 151872 5438
rect 151820 5374 151872 5380
rect 150624 3324 150676 3330
rect 150624 3266 150676 3272
rect 151728 3324 151780 3330
rect 151728 3266 151780 3272
rect 150636 480 150664 3266
rect 151832 480 151860 5374
rect 153028 480 153056 5782
rect 153212 3262 153240 60030
rect 155972 57186 156000 60044
rect 158548 57934 158576 60044
rect 158536 57928 158588 57934
rect 158536 57870 158588 57876
rect 155960 57180 156012 57186
rect 155960 57122 156012 57128
rect 157340 56976 157392 56982
rect 157340 56918 157392 56924
rect 160008 56976 160060 56982
rect 160008 56918 160060 56924
rect 155866 17504 155922 17513
rect 155866 17439 155922 17448
rect 154210 7712 154266 7721
rect 154210 7647 154266 7656
rect 153200 3256 153252 3262
rect 153200 3198 153252 3204
rect 154224 480 154252 7647
rect 155880 3330 155908 17439
rect 157352 16574 157380 56918
rect 157352 16546 157840 16574
rect 156604 4888 156656 4894
rect 156604 4830 156656 4836
rect 155408 3324 155460 3330
rect 155408 3266 155460 3272
rect 155868 3324 155920 3330
rect 155868 3266 155920 3272
rect 155420 480 155448 3266
rect 156616 480 156644 4830
rect 157812 480 157840 16546
rect 160020 3330 160048 56918
rect 160112 4214 160140 60522
rect 161138 60030 161428 60058
rect 160192 8288 160244 8294
rect 160192 8230 160244 8236
rect 160100 4208 160152 4214
rect 160100 4150 160152 4156
rect 160204 3482 160232 8230
rect 161400 4894 161428 60030
rect 164148 56840 164200 56846
rect 164148 56782 164200 56788
rect 162766 21448 162822 21457
rect 162766 21383 162822 21392
rect 162780 6914 162808 21383
rect 162504 6886 162808 6914
rect 161388 4888 161440 4894
rect 161388 4830 161440 4836
rect 161296 4208 161348 4214
rect 161296 4150 161348 4156
rect 160112 3454 160232 3482
rect 158904 3324 158956 3330
rect 158904 3266 158956 3272
rect 160008 3324 160060 3330
rect 160008 3266 160060 3272
rect 158916 480 158944 3266
rect 160112 480 160140 3454
rect 161308 480 161336 4150
rect 162504 480 162532 6886
rect 164160 3330 164188 56782
rect 164344 56778 164372 60044
rect 164332 56772 164384 56778
rect 164332 56714 164384 56720
rect 166920 47598 166948 60044
rect 166908 47592 166960 47598
rect 166908 47534 166960 47540
rect 166908 13388 166960 13394
rect 166908 13330 166960 13336
rect 164884 5228 164936 5234
rect 164884 5170 164936 5176
rect 163688 3324 163740 3330
rect 163688 3266 163740 3272
rect 164148 3324 164200 3330
rect 164148 3266 164200 3272
rect 163700 480 163728 3266
rect 164896 480 164924 5170
rect 166920 3330 166948 13330
rect 166080 3324 166132 3330
rect 166080 3266 166132 3272
rect 166908 3324 166960 3330
rect 166908 3266 166960 3272
rect 166092 480 166120 3266
rect 168300 3262 168328 60522
rect 169510 60030 169708 60058
rect 168380 59900 168432 59906
rect 168380 59842 168432 59848
rect 167184 3256 167236 3262
rect 167184 3198 167236 3204
rect 168288 3256 168340 3262
rect 168288 3198 168340 3204
rect 167196 480 167224 3198
rect 168392 480 168420 59842
rect 169576 8288 169628 8294
rect 169576 8230 169628 8236
rect 169588 480 169616 8230
rect 169680 4418 169708 60030
rect 171048 58948 171100 58954
rect 171048 58890 171100 58896
rect 171060 6914 171088 58890
rect 172716 57934 172744 60044
rect 173900 59968 173952 59974
rect 173900 59910 173952 59916
rect 172704 57928 172756 57934
rect 172704 57870 172756 57876
rect 173808 57928 173860 57934
rect 173808 57870 173860 57876
rect 173820 15978 173848 57870
rect 173912 16574 173940 59910
rect 175292 57186 175320 60044
rect 175280 57180 175332 57186
rect 175280 57122 175332 57128
rect 173912 16546 174308 16574
rect 173808 15972 173860 15978
rect 173808 15914 173860 15920
rect 173164 7540 173216 7546
rect 173164 7482 173216 7488
rect 170784 6886 171088 6914
rect 169668 4412 169720 4418
rect 169668 4354 169720 4360
rect 170784 480 170812 6886
rect 171968 5228 172020 5234
rect 171968 5170 172020 5176
rect 171980 480 172008 5170
rect 173176 480 173204 7482
rect 174280 480 174308 16546
rect 176568 14612 176620 14618
rect 176568 14554 176620 14560
rect 176580 3330 176608 14554
rect 176672 3330 176700 60590
rect 177882 60030 177988 60058
rect 177960 6798 177988 60030
rect 180444 57934 180472 60044
rect 180432 57928 180484 57934
rect 180432 57870 180484 57876
rect 182088 57044 182140 57050
rect 182088 56986 182140 56992
rect 178040 56432 178092 56438
rect 178040 56374 178092 56380
rect 178052 16574 178080 56374
rect 180708 54868 180760 54874
rect 180708 54810 180760 54816
rect 178052 16546 179092 16574
rect 176752 6792 176804 6798
rect 176752 6734 176804 6740
rect 177948 6792 178000 6798
rect 177948 6734 178000 6740
rect 175464 3324 175516 3330
rect 175464 3266 175516 3272
rect 176568 3324 176620 3330
rect 176568 3266 176620 3272
rect 176660 3324 176712 3330
rect 176660 3266 176712 3272
rect 175476 480 175504 3266
rect 176764 3210 176792 6734
rect 177856 3324 177908 3330
rect 177856 3266 177908 3272
rect 176672 3182 176792 3210
rect 176672 480 176700 3182
rect 177868 480 177896 3266
rect 179064 480 179092 16546
rect 180720 3330 180748 54810
rect 182100 3330 182128 56986
rect 183664 56778 183692 60044
rect 186240 58410 186268 60044
rect 186228 58404 186280 58410
rect 186228 58346 186280 58352
rect 188816 57934 188844 60044
rect 188988 58608 189040 58614
rect 188988 58550 189040 58556
rect 184940 57928 184992 57934
rect 184940 57870 184992 57876
rect 188804 57928 188856 57934
rect 188804 57870 188856 57876
rect 183652 56772 183704 56778
rect 183652 56714 183704 56720
rect 184848 53440 184900 53446
rect 184848 53382 184900 53388
rect 183468 11892 183520 11898
rect 183468 11834 183520 11840
rect 183480 3330 183508 11834
rect 180248 3324 180300 3330
rect 180248 3266 180300 3272
rect 180708 3324 180760 3330
rect 180708 3266 180760 3272
rect 181444 3324 181496 3330
rect 181444 3266 181496 3272
rect 182088 3324 182140 3330
rect 182088 3266 182140 3272
rect 182548 3324 182600 3330
rect 182548 3266 182600 3272
rect 183468 3324 183520 3330
rect 183468 3266 183520 3272
rect 180260 480 180288 3266
rect 181456 480 181484 3266
rect 182560 480 182588 3266
rect 184860 3262 184888 53382
rect 183744 3256 183796 3262
rect 183744 3198 183796 3204
rect 184848 3256 184900 3262
rect 184848 3198 184900 3204
rect 183756 480 183784 3198
rect 184952 480 184980 57870
rect 186136 11960 186188 11966
rect 186136 11902 186188 11908
rect 186148 480 186176 11902
rect 187332 6588 187384 6594
rect 187332 6530 187384 6536
rect 187344 480 187372 6530
rect 189000 3330 189028 58550
rect 191392 58342 191420 60044
rect 191380 58336 191432 58342
rect 191380 58278 191432 58284
rect 194612 57730 194640 60044
rect 191840 57724 191892 57730
rect 191840 57666 191892 57672
rect 194600 57724 194652 57730
rect 194600 57666 194652 57672
rect 195888 57724 195940 57730
rect 195888 57666 195940 57672
rect 191748 56432 191800 56438
rect 191748 56374 191800 56380
rect 190368 11960 190420 11966
rect 190368 11902 190420 11908
rect 190380 3330 190408 11902
rect 191760 3330 191788 56374
rect 191852 16574 191880 57666
rect 194692 56772 194744 56778
rect 194692 56714 194744 56720
rect 194704 45554 194732 56714
rect 194612 45526 194732 45554
rect 194612 16574 194640 45526
rect 191852 16546 192064 16574
rect 194612 16546 195652 16574
rect 188528 3324 188580 3330
rect 188528 3266 188580 3272
rect 188988 3324 189040 3330
rect 188988 3266 189040 3272
rect 189724 3324 189776 3330
rect 189724 3266 189776 3272
rect 190368 3324 190420 3330
rect 190368 3266 190420 3272
rect 190828 3324 190880 3330
rect 190828 3266 190880 3272
rect 191748 3324 191800 3330
rect 191748 3266 191800 3272
rect 188540 480 188568 3266
rect 189736 480 189764 3266
rect 190840 480 190868 3266
rect 192036 480 192064 16546
rect 194416 8152 194468 8158
rect 194416 8094 194468 8100
rect 193218 4176 193274 4185
rect 193218 4111 193274 4120
rect 193232 480 193260 4111
rect 194428 480 194456 8094
rect 195624 480 195652 16546
rect 195900 6594 195928 57666
rect 197188 56914 197216 60044
rect 199778 60030 199976 60058
rect 197176 56908 197228 56914
rect 197176 56850 197228 56856
rect 197912 9444 197964 9450
rect 197912 9386 197964 9392
rect 195888 6588 195940 6594
rect 195888 6530 195940 6536
rect 196808 5296 196860 5302
rect 196808 5238 196860 5244
rect 196820 480 196848 5238
rect 197924 480 197952 9386
rect 199948 7070 199976 60030
rect 199936 7064 199988 7070
rect 199936 7006 199988 7012
rect 200040 3330 200068 60590
rect 336740 60512 336792 60518
rect 336740 60454 336792 60460
rect 350448 60512 350500 60518
rect 350448 60454 350500 60460
rect 358728 60512 358780 60518
rect 358728 60454 358780 60460
rect 202788 59968 202840 59974
rect 202788 59910 202840 59916
rect 201500 58472 201552 58478
rect 201500 58414 201552 58420
rect 200120 56500 200172 56506
rect 200120 56442 200172 56448
rect 200132 16574 200160 56442
rect 200132 16546 200344 16574
rect 199108 3324 199160 3330
rect 199108 3266 199160 3272
rect 200028 3324 200080 3330
rect 200028 3266 200080 3272
rect 199120 480 199148 3266
rect 200316 480 200344 16546
rect 201512 480 201540 58414
rect 202800 6914 202828 59910
rect 202984 57526 203012 60044
rect 204272 60030 205574 60058
rect 208150 60030 208348 60058
rect 202972 57520 203024 57526
rect 202972 57462 203024 57468
rect 203892 7200 203944 7206
rect 203892 7142 203944 7148
rect 202708 6886 202828 6914
rect 202708 480 202736 6886
rect 203904 480 203932 7142
rect 204272 4486 204300 60030
rect 205640 57112 205692 57118
rect 205640 57054 205692 57060
rect 205652 16574 205680 57054
rect 205652 16546 206232 16574
rect 205546 11792 205602 11801
rect 205546 11727 205602 11736
rect 204260 4480 204312 4486
rect 204260 4422 204312 4428
rect 205560 3330 205588 11727
rect 205088 3324 205140 3330
rect 205088 3266 205140 3272
rect 205548 3324 205600 3330
rect 205548 3266 205600 3272
rect 205100 480 205128 3266
rect 206204 480 206232 16546
rect 208216 12028 208268 12034
rect 208216 11970 208268 11976
rect 208228 3330 208256 11970
rect 208320 5302 208348 60030
rect 210712 57730 210740 60044
rect 211068 59900 211120 59906
rect 211068 59842 211120 59848
rect 209872 57724 209924 57730
rect 209872 57666 209924 57672
rect 210700 57724 210752 57730
rect 210700 57666 210752 57672
rect 209780 53508 209832 53514
rect 209780 53450 209832 53456
rect 209688 22840 209740 22846
rect 209688 22782 209740 22788
rect 208308 5296 208360 5302
rect 208308 5238 208360 5244
rect 209700 3330 209728 22782
rect 207388 3324 207440 3330
rect 207388 3266 207440 3272
rect 208216 3324 208268 3330
rect 208216 3266 208268 3272
rect 208584 3324 208636 3330
rect 208584 3266 208636 3272
rect 209688 3324 209740 3330
rect 209688 3266 209740 3272
rect 207400 480 207428 3266
rect 208596 480 208624 3266
rect 209792 480 209820 53450
rect 209884 51814 209912 57666
rect 209872 51808 209924 51814
rect 209872 51750 209924 51756
rect 211080 6914 211108 59842
rect 213828 57724 213880 57730
rect 213828 57666 213880 57672
rect 212448 56908 212500 56914
rect 212448 56850 212500 56856
rect 212460 6914 212488 56850
rect 210988 6886 211108 6914
rect 212184 6886 212488 6914
rect 210988 480 211016 6886
rect 212184 480 212212 6886
rect 213840 3398 213868 57666
rect 213932 52086 213960 60044
rect 216522 60030 216628 60058
rect 219098 60030 219388 60058
rect 213920 52080 213972 52086
rect 213920 52022 213972 52028
rect 216600 16046 216628 60030
rect 218060 59900 218112 59906
rect 218060 59842 218112 59848
rect 217966 18728 218022 18737
rect 217966 18663 218022 18672
rect 214472 16040 214524 16046
rect 214472 15982 214524 15988
rect 216588 16040 216640 16046
rect 216588 15982 216640 15988
rect 213368 3392 213420 3398
rect 213368 3334 213420 3340
rect 213828 3392 213880 3398
rect 213828 3334 213880 3340
rect 213380 480 213408 3334
rect 214484 480 214512 15982
rect 216586 12064 216642 12073
rect 216586 11999 216642 12008
rect 216600 3398 216628 11999
rect 217980 3398 218008 18663
rect 218072 16574 218100 59842
rect 218072 16546 219204 16574
rect 219176 3482 219204 16546
rect 219256 13320 219308 13326
rect 219256 13262 219308 13268
rect 219268 6914 219296 13262
rect 219360 8158 219388 60030
rect 220832 60030 221674 60058
rect 224788 60030 224894 60058
rect 227470 60030 227576 60058
rect 220728 57112 220780 57118
rect 220728 57054 220780 57060
rect 219348 8152 219400 8158
rect 219348 8094 219400 8100
rect 220740 6914 220768 57054
rect 219268 6886 219388 6914
rect 219176 3454 219296 3482
rect 215668 3392 215720 3398
rect 215668 3334 215720 3340
rect 216588 3392 216640 3398
rect 216588 3334 216640 3340
rect 216864 3392 216916 3398
rect 216864 3334 216916 3340
rect 217968 3392 218020 3398
rect 217968 3334 218020 3340
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 215680 480 215708 3334
rect 216876 480 216904 3334
rect 218072 480 218100 3334
rect 219268 480 219296 3454
rect 219360 3398 219388 6886
rect 220464 6886 220768 6914
rect 219348 3392 219400 3398
rect 219348 3334 219400 3340
rect 220464 480 220492 6886
rect 220832 3330 220860 60030
rect 224684 59900 224736 59906
rect 224684 59842 224736 59848
rect 220912 28280 220964 28286
rect 220912 28222 220964 28228
rect 220924 16574 220952 28222
rect 220924 16546 221596 16574
rect 220820 3324 220872 3330
rect 220820 3266 220872 3272
rect 221568 480 221596 16546
rect 222752 9648 222804 9654
rect 222752 9590 222804 9596
rect 222764 480 222792 9590
rect 224696 3398 224724 59842
rect 224788 7274 224816 60030
rect 226524 57860 226576 57866
rect 226524 57802 226576 57808
rect 224776 7268 224828 7274
rect 224776 7210 224828 7216
rect 226536 6914 226564 57802
rect 227548 7478 227576 60030
rect 227628 59900 227680 59906
rect 227628 59842 227680 59848
rect 227536 7472 227588 7478
rect 227536 7414 227588 7420
rect 227640 6914 227668 59842
rect 229192 59832 229244 59838
rect 229192 59774 229244 59780
rect 229204 16574 229232 59774
rect 230032 56846 230060 60044
rect 233148 58472 233200 58478
rect 233148 58414 233200 58420
rect 230020 56840 230072 56846
rect 230020 56782 230072 56788
rect 229204 16546 229876 16574
rect 228732 7132 228784 7138
rect 228732 7074 228784 7080
rect 226352 6886 226564 6914
rect 227548 6886 227668 6914
rect 225144 5432 225196 5438
rect 225144 5374 225196 5380
rect 223948 3392 224000 3398
rect 223948 3334 224000 3340
rect 224684 3392 224736 3398
rect 224684 3334 224736 3340
rect 223960 480 223988 3334
rect 225156 480 225184 5374
rect 226352 480 226380 6886
rect 227548 480 227576 6886
rect 228744 480 228772 7074
rect 229848 480 229876 16546
rect 231766 14648 231822 14657
rect 231766 14583 231822 14592
rect 231780 3398 231808 14583
rect 233160 3398 233188 58414
rect 233252 57526 233280 60044
rect 234632 60030 235842 60058
rect 234528 57860 234580 57866
rect 234528 57802 234580 57808
rect 233240 57520 233292 57526
rect 233240 57462 233292 57468
rect 234436 57520 234488 57526
rect 234436 57462 234488 57468
rect 234448 4350 234476 57462
rect 234436 4344 234488 4350
rect 234436 4286 234488 4292
rect 234540 3398 234568 57802
rect 234632 4962 234660 60030
rect 236000 59832 236052 59838
rect 236000 59774 236052 59780
rect 236012 16574 236040 59774
rect 238404 59090 238432 60044
rect 238392 59084 238444 59090
rect 238392 59026 238444 59032
rect 240980 57526 241008 60044
rect 240968 57520 241020 57526
rect 240968 57462 241020 57468
rect 237378 26888 237434 26897
rect 237378 26823 237434 26832
rect 237392 16574 237420 26823
rect 236012 16546 237052 16574
rect 237392 16546 238156 16574
rect 234712 7336 234764 7342
rect 234712 7278 234764 7284
rect 234620 4956 234672 4962
rect 234620 4898 234672 4904
rect 234724 3482 234752 7278
rect 235814 4176 235870 4185
rect 235814 4111 235870 4120
rect 234632 3454 234752 3482
rect 231032 3392 231084 3398
rect 231032 3334 231084 3340
rect 231768 3392 231820 3398
rect 231768 3334 231820 3340
rect 232228 3392 232280 3398
rect 232228 3334 232280 3340
rect 233148 3392 233200 3398
rect 233148 3334 233200 3340
rect 233424 3392 233476 3398
rect 233424 3334 233476 3340
rect 234528 3392 234580 3398
rect 234528 3334 234580 3340
rect 231044 480 231072 3334
rect 232240 480 232268 3334
rect 233436 480 233464 3334
rect 234632 480 234660 3454
rect 235828 480 235856 4111
rect 237024 480 237052 16546
rect 238128 480 238156 16546
rect 240506 14512 240562 14521
rect 240506 14447 240562 14456
rect 239312 4480 239364 4486
rect 239312 4422 239364 4428
rect 239324 480 239352 4422
rect 240520 480 240548 14447
rect 241704 7064 241756 7070
rect 241704 7006 241756 7012
rect 241716 480 241744 7006
rect 244094 5672 244150 5681
rect 244094 5607 244150 5616
rect 242900 4344 242952 4350
rect 242900 4286 242952 4292
rect 242912 480 242940 4286
rect 244108 480 244136 5607
rect 244200 4962 244228 60044
rect 245672 60030 246790 60058
rect 244280 57452 244332 57458
rect 244280 57394 244332 57400
rect 244292 16574 244320 57394
rect 245672 45558 245700 60030
rect 248328 59832 248380 59838
rect 248328 59774 248380 59780
rect 245660 45552 245712 45558
rect 245660 45494 245712 45500
rect 244292 16546 245240 16574
rect 244188 4956 244240 4962
rect 244188 4898 244240 4904
rect 245212 480 245240 16546
rect 246394 15872 246450 15881
rect 246394 15807 246450 15816
rect 246408 480 246436 15807
rect 248340 3398 248368 59774
rect 249352 56982 249380 60044
rect 249340 56976 249392 56982
rect 249340 56918 249392 56924
rect 251928 56914 251956 60044
rect 254032 59764 254084 59770
rect 254032 59706 254084 59712
rect 251916 56908 251968 56914
rect 251916 56850 251968 56856
rect 249708 55072 249760 55078
rect 249708 55014 249760 55020
rect 249720 3398 249748 55014
rect 252466 24168 252522 24177
rect 252466 24103 252522 24112
rect 252376 8696 252428 8702
rect 252376 8638 252428 8644
rect 249984 4684 250036 4690
rect 249984 4626 250036 4632
rect 247592 3392 247644 3398
rect 247592 3334 247644 3340
rect 248328 3392 248380 3398
rect 248328 3334 248380 3340
rect 248788 3392 248840 3398
rect 248788 3334 248840 3340
rect 249708 3392 249760 3398
rect 249708 3334 249760 3340
rect 247604 480 247632 3334
rect 248800 480 248828 3334
rect 249996 480 250024 4626
rect 251180 3392 251232 3398
rect 251180 3334 251232 3340
rect 251192 480 251220 3334
rect 252388 480 252416 8638
rect 252480 3398 252508 24103
rect 254044 16574 254072 59706
rect 255148 57866 255176 60044
rect 257738 60030 257936 60058
rect 260314 60030 260788 60058
rect 262890 60030 263548 60058
rect 266110 60030 266308 60058
rect 268686 60030 269068 60058
rect 255136 57860 255188 57866
rect 255136 57802 255188 57808
rect 255320 55004 255372 55010
rect 255320 54946 255372 54952
rect 255332 16574 255360 54946
rect 254044 16546 254716 16574
rect 255332 16546 255912 16574
rect 253478 10976 253534 10985
rect 253478 10911 253534 10920
rect 252468 3392 252520 3398
rect 252468 3334 252520 3340
rect 253492 480 253520 10911
rect 254688 480 254716 16546
rect 255884 480 255912 16546
rect 257908 7002 257936 60030
rect 257988 59764 258040 59770
rect 257988 59706 258040 59712
rect 258080 59764 258132 59770
rect 258080 59706 258132 59712
rect 257896 6996 257948 7002
rect 257896 6938 257948 6944
rect 258000 3398 258028 59706
rect 258092 16574 258120 59706
rect 258092 16546 258304 16574
rect 257068 3392 257120 3398
rect 257068 3334 257120 3340
rect 257988 3392 258040 3398
rect 257988 3334 258040 3340
rect 257080 480 257108 3334
rect 258276 480 258304 16546
rect 260760 14754 260788 60030
rect 260748 14748 260800 14754
rect 260748 14690 260800 14696
rect 262956 8628 263008 8634
rect 262956 8570 263008 8576
rect 259460 8492 259512 8498
rect 259460 8434 259512 8440
rect 259472 480 259500 8434
rect 261758 5672 261814 5681
rect 261758 5607 261814 5616
rect 260656 4684 260708 4690
rect 260656 4626 260708 4632
rect 260668 480 260696 4626
rect 261772 480 261800 5607
rect 262968 480 262996 8570
rect 263520 7342 263548 60030
rect 265348 8560 265400 8566
rect 265348 8502 265400 8508
rect 263508 7336 263560 7342
rect 263508 7278 263560 7284
rect 264152 4752 264204 4758
rect 264152 4694 264204 4700
rect 264164 480 264192 4694
rect 265360 480 265388 8502
rect 266280 7070 266308 60030
rect 269040 14686 269068 60030
rect 271248 59090 271276 60044
rect 273272 60030 274482 60058
rect 277058 60030 277348 60058
rect 271236 59084 271288 59090
rect 271236 59026 271288 59032
rect 273168 57452 273220 57458
rect 273168 57394 273220 57400
rect 269028 14680 269080 14686
rect 269028 14622 269080 14628
rect 270040 8900 270092 8906
rect 270040 8842 270092 8848
rect 266544 8832 266596 8838
rect 266544 8774 266596 8780
rect 266268 7064 266320 7070
rect 266268 7006 266320 7012
rect 266556 480 266584 8774
rect 268844 8764 268896 8770
rect 268844 8706 268896 8712
rect 267740 4616 267792 4622
rect 267740 4558 267792 4564
rect 267752 480 267780 4558
rect 268856 480 268884 8706
rect 270052 480 270080 8842
rect 271236 4412 271288 4418
rect 271236 4354 271288 4360
rect 271248 480 271276 4354
rect 273180 3398 273208 57394
rect 273272 6118 273300 60030
rect 274548 56500 274600 56506
rect 274548 56442 274600 56448
rect 273260 6112 273312 6118
rect 273260 6054 273312 6060
rect 274560 3398 274588 56442
rect 277320 28286 277348 60030
rect 279620 57594 279648 60044
rect 282196 57866 282224 60044
rect 282184 57860 282236 57866
rect 282184 57802 282236 57808
rect 284208 57860 284260 57866
rect 284208 57802 284260 57808
rect 279608 57588 279660 57594
rect 279608 57530 279660 57536
rect 282184 57588 282236 57594
rect 282184 57530 282236 57536
rect 277308 28280 277360 28286
rect 277308 28222 277360 28228
rect 281538 17368 281594 17377
rect 281538 17303 281594 17312
rect 281552 16574 281580 17303
rect 282196 17270 282224 57530
rect 282184 17264 282236 17270
rect 282184 17206 282236 17212
rect 281552 16546 281948 16574
rect 277124 9580 277176 9586
rect 277124 9522 277176 9528
rect 274824 4752 274876 4758
rect 274824 4694 274876 4700
rect 272432 3392 272484 3398
rect 272432 3334 272484 3340
rect 273168 3392 273220 3398
rect 273168 3334 273220 3340
rect 273628 3392 273680 3398
rect 273628 3334 273680 3340
rect 274548 3392 274600 3398
rect 274548 3334 274600 3340
rect 272444 480 272472 3334
rect 273640 480 273668 3334
rect 274836 480 274864 4694
rect 276018 4176 276074 4185
rect 276018 4111 276074 4120
rect 276032 480 276060 4111
rect 277136 480 277164 9522
rect 280712 9512 280764 9518
rect 280712 9454 280764 9460
rect 278320 4616 278372 4622
rect 278320 4558 278372 4564
rect 278332 480 278360 4558
rect 279514 4176 279570 4185
rect 279514 4111 279570 4120
rect 279528 480 279556 4111
rect 280724 480 280752 9454
rect 281920 480 281948 16546
rect 284220 3398 284248 57802
rect 285416 57050 285444 60044
rect 286968 59764 287020 59770
rect 286968 59706 287020 59712
rect 285404 57044 285456 57050
rect 285404 56986 285456 56992
rect 284300 54936 284352 54942
rect 284300 54878 284352 54884
rect 284312 16574 284340 54878
rect 285588 53508 285640 53514
rect 285588 53450 285640 53456
rect 284312 16546 285444 16574
rect 283104 3392 283156 3398
rect 283104 3334 283156 3340
rect 284208 3392 284260 3398
rect 284208 3334 284260 3340
rect 284300 3392 284352 3398
rect 284300 3334 284352 3340
rect 283116 480 283144 3334
rect 284312 480 284340 3334
rect 285416 480 285444 16546
rect 285600 3398 285628 53450
rect 286980 6914 287008 59706
rect 287992 57798 288020 60044
rect 289832 60030 290582 60058
rect 287980 57792 288032 57798
rect 287980 57734 288032 57740
rect 287060 57656 287112 57662
rect 287060 57598 287112 57604
rect 287072 16574 287100 57598
rect 288440 52012 288492 52018
rect 288440 51954 288492 51960
rect 288452 16574 288480 51954
rect 287072 16546 287836 16574
rect 288452 16546 289032 16574
rect 286612 6886 287008 6914
rect 285588 3392 285640 3398
rect 285588 3334 285640 3340
rect 286612 480 286640 6886
rect 287808 480 287836 16546
rect 289004 480 289032 16546
rect 289832 5914 289860 60030
rect 291108 59764 291160 59770
rect 291108 59706 291160 59712
rect 289820 5908 289872 5914
rect 289820 5850 289872 5856
rect 291120 3398 291148 59706
rect 293144 59022 293172 60044
rect 293132 59016 293184 59022
rect 293132 58958 293184 58964
rect 296364 57458 296392 60044
rect 296720 58540 296772 58546
rect 296720 58482 296772 58488
rect 296352 57452 296404 57458
rect 296352 57394 296404 57400
rect 291200 57180 291252 57186
rect 291200 57122 291252 57128
rect 291212 16574 291240 57122
rect 295984 56636 296036 56642
rect 295984 56578 296036 56584
rect 295248 53576 295300 53582
rect 295248 53518 295300 53524
rect 291212 16546 291424 16574
rect 290188 3392 290240 3398
rect 290188 3334 290240 3340
rect 291108 3392 291160 3398
rect 291108 3334 291160 3340
rect 290200 480 290228 3334
rect 291396 480 291424 16546
rect 293682 10432 293738 10441
rect 293682 10367 293738 10376
rect 292580 4344 292632 4350
rect 292580 4286 292632 4292
rect 292592 480 292620 4286
rect 293696 480 293724 10367
rect 295260 6914 295288 53518
rect 295996 13394 296024 56578
rect 296732 16574 296760 58482
rect 298744 57520 298796 57526
rect 298744 57462 298796 57468
rect 296732 16546 297312 16574
rect 296626 15872 296682 15881
rect 296626 15807 296682 15816
rect 295984 13388 296036 13394
rect 295984 13330 296036 13336
rect 294892 6886 295288 6914
rect 294892 480 294920 6886
rect 296640 3398 296668 15807
rect 296076 3392 296128 3398
rect 296076 3334 296128 3340
rect 296628 3392 296680 3398
rect 296628 3334 296680 3340
rect 296088 480 296116 3334
rect 297284 480 297312 16546
rect 298756 4418 298784 57462
rect 298940 56642 298968 60044
rect 301516 57458 301544 60044
rect 302240 59764 302292 59770
rect 302240 59706 302292 59712
rect 301504 57452 301556 57458
rect 301504 57394 301556 57400
rect 299480 57384 299532 57390
rect 299480 57326 299532 57332
rect 298928 56636 298980 56642
rect 298928 56578 298980 56584
rect 299388 26920 299440 26926
rect 299388 26862 299440 26868
rect 298744 4412 298796 4418
rect 298744 4354 298796 4360
rect 299400 3398 299428 26862
rect 299492 3398 299520 57326
rect 302252 16574 302280 59706
rect 304736 57390 304764 60044
rect 306392 60030 307326 60058
rect 304724 57384 304776 57390
rect 304724 57326 304776 57332
rect 302252 16546 303200 16574
rect 301964 6112 302016 6118
rect 301964 6054 302016 6060
rect 299664 4548 299716 4554
rect 299664 4490 299716 4496
rect 298468 3392 298520 3398
rect 298468 3334 298520 3340
rect 299388 3392 299440 3398
rect 299388 3334 299440 3340
rect 299480 3392 299532 3398
rect 299480 3334 299532 3340
rect 298480 480 298508 3334
rect 299676 480 299704 4490
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 300780 480 300808 3334
rect 301976 480 302004 6054
rect 303172 480 303200 16546
rect 304356 9376 304408 9382
rect 304356 9318 304408 9324
rect 304368 480 304396 9318
rect 306392 5982 306420 60030
rect 307760 57928 307812 57934
rect 307760 57870 307812 57876
rect 306380 5976 306432 5982
rect 306380 5918 306432 5924
rect 306748 5364 306800 5370
rect 306748 5306 306800 5312
rect 305550 3088 305606 3097
rect 305550 3023 305606 3032
rect 305564 480 305592 3023
rect 306760 480 306788 5306
rect 307772 3482 307800 57870
rect 309888 57526 309916 60044
rect 311912 60030 312478 60058
rect 314672 60030 315698 60058
rect 317432 60030 318274 60058
rect 309876 57520 309928 57526
rect 309876 57462 309928 57468
rect 310428 52012 310480 52018
rect 310428 51954 310480 51960
rect 307850 11928 307906 11937
rect 307850 11863 307906 11872
rect 307864 3874 307892 11863
rect 310440 6914 310468 51954
rect 311440 9308 311492 9314
rect 311440 9250 311492 9256
rect 310256 6886 310468 6914
rect 307852 3868 307904 3874
rect 307852 3810 307904 3816
rect 309048 3868 309100 3874
rect 309048 3810 309100 3816
rect 307772 3454 307984 3482
rect 307956 480 307984 3454
rect 309060 480 309088 3810
rect 310256 480 310284 6886
rect 311452 480 311480 9250
rect 311912 4010 311940 60030
rect 312636 9240 312688 9246
rect 312636 9182 312688 9188
rect 311900 4004 311952 4010
rect 311900 3946 311952 3952
rect 312648 480 312676 9182
rect 313832 4548 313884 4554
rect 313832 4490 313884 4496
rect 313844 480 313872 4490
rect 314672 3398 314700 60030
rect 315948 59764 316000 59770
rect 315948 59706 316000 59712
rect 315960 3398 315988 59706
rect 317432 6050 317460 60030
rect 320836 59158 320864 60044
rect 320824 59152 320876 59158
rect 320824 59094 320876 59100
rect 323412 57662 323440 60044
rect 326632 57798 326660 60044
rect 326620 57792 326672 57798
rect 326620 57734 326672 57740
rect 323400 57656 323452 57662
rect 323400 57598 323452 57604
rect 324228 57656 324280 57662
rect 324228 57598 324280 57604
rect 320824 57520 320876 57526
rect 320824 57462 320876 57468
rect 319720 10804 319772 10810
rect 319720 10746 319772 10752
rect 318524 9172 318576 9178
rect 318524 9114 318576 9120
rect 317420 6044 317472 6050
rect 317420 5986 317472 5992
rect 317328 5500 317380 5506
rect 317328 5442 317380 5448
rect 316224 5364 316276 5370
rect 316224 5306 316276 5312
rect 314660 3392 314712 3398
rect 314660 3334 314712 3340
rect 315028 3392 315080 3398
rect 315028 3334 315080 3340
rect 315948 3392 316000 3398
rect 315948 3334 316000 3340
rect 315040 480 315068 3334
rect 316236 480 316264 5306
rect 317340 480 317368 5442
rect 318536 480 318564 9114
rect 319732 480 319760 10746
rect 320836 9178 320864 57462
rect 322938 17232 322994 17241
rect 322938 17167 322994 17176
rect 322952 16574 322980 17167
rect 322952 16546 323348 16574
rect 320824 9172 320876 9178
rect 320824 9114 320876 9120
rect 320916 6996 320968 7002
rect 320916 6938 320968 6944
rect 320928 480 320956 6938
rect 322112 6044 322164 6050
rect 322112 5986 322164 5992
rect 322124 480 322152 5986
rect 323320 480 323348 16546
rect 324240 6914 324268 57598
rect 329208 57526 329236 60044
rect 329196 57520 329248 57526
rect 329196 57462 329248 57468
rect 331784 57118 331812 60044
rect 335018 60030 335308 60058
rect 331772 57112 331824 57118
rect 331772 57054 331824 57060
rect 324320 56364 324372 56370
rect 324320 56306 324372 56312
rect 324148 6886 324268 6914
rect 324148 3874 324176 6886
rect 324136 3868 324188 3874
rect 324136 3810 324188 3816
rect 324332 3398 324360 56306
rect 325700 22772 325752 22778
rect 325700 22714 325752 22720
rect 325712 16574 325740 22714
rect 335280 17270 335308 60030
rect 328460 17264 328512 17270
rect 328460 17206 328512 17212
rect 335268 17264 335320 17270
rect 335268 17206 335320 17212
rect 328472 16574 328500 17206
rect 325712 16546 326844 16574
rect 328472 16546 329236 16574
rect 324412 5092 324464 5098
rect 324412 5034 324464 5040
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 324424 480 324452 5034
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 326816 480 326844 16546
rect 328000 4276 328052 4282
rect 328000 4218 328052 4224
rect 328012 480 328040 4218
rect 329208 480 329236 16546
rect 332506 15872 332562 15881
rect 332506 15807 332562 15816
rect 330392 5976 330444 5982
rect 330392 5918 330444 5924
rect 329838 3088 329894 3097
rect 329838 3023 329840 3032
rect 329892 3023 329894 3032
rect 329840 2994 329892 3000
rect 330404 480 330432 5918
rect 332520 3398 332548 15807
rect 336278 9616 336334 9625
rect 336278 9551 336334 9560
rect 332690 5672 332746 5681
rect 332690 5607 332746 5616
rect 331588 3392 331640 3398
rect 331588 3334 331640 3340
rect 332508 3392 332560 3398
rect 332508 3334 332560 3340
rect 331600 480 331628 3334
rect 332704 480 332732 5607
rect 335084 5092 335136 5098
rect 335084 5034 335136 5040
rect 333886 4176 333942 4185
rect 333886 4111 333942 4120
rect 333900 480 333928 4111
rect 335096 480 335124 5034
rect 336292 480 336320 9551
rect 336752 6914 336780 60454
rect 336844 60030 337594 60058
rect 339512 60030 340170 60058
rect 336844 7206 336872 60030
rect 338120 53372 338172 53378
rect 338120 53314 338172 53320
rect 338132 16574 338160 53314
rect 338132 16546 338712 16574
rect 336832 7200 336884 7206
rect 336832 7142 336884 7148
rect 336752 6886 337516 6914
rect 337488 480 337516 6886
rect 338684 480 338712 16546
rect 339512 4350 339540 60030
rect 342732 59158 342760 60044
rect 342720 59152 342772 59158
rect 342720 59094 342772 59100
rect 345952 58546 345980 60044
rect 347792 60030 348542 60058
rect 345940 58540 345992 58546
rect 345940 58482 345992 58488
rect 343548 57656 343600 57662
rect 343548 57598 343600 57604
rect 342166 40624 342222 40633
rect 342166 40559 342222 40568
rect 339868 15904 339920 15910
rect 339868 15846 339920 15852
rect 339500 4344 339552 4350
rect 339500 4286 339552 4292
rect 339880 480 339908 15846
rect 342076 7404 342128 7410
rect 342076 7346 342128 7352
rect 340972 4004 341024 4010
rect 340972 3946 341024 3952
rect 340984 480 341012 3946
rect 342088 3482 342116 7346
rect 342180 4010 342208 40559
rect 343560 6914 343588 57598
rect 346308 56364 346360 56370
rect 346308 56306 346360 56312
rect 344558 8936 344614 8945
rect 344558 8871 344614 8880
rect 343376 6886 343588 6914
rect 342168 4004 342220 4010
rect 342168 3946 342220 3952
rect 342088 3454 342208 3482
rect 342180 480 342208 3454
rect 343376 480 343404 6886
rect 344572 480 344600 8871
rect 346320 3398 346348 56306
rect 346952 9104 347004 9110
rect 346952 9046 347004 9052
rect 345756 3392 345808 3398
rect 345756 3334 345808 3340
rect 346308 3392 346360 3398
rect 346308 3334 346360 3340
rect 345768 480 345796 3334
rect 346964 480 346992 9046
rect 347792 3942 347820 60030
rect 349160 54800 349212 54806
rect 349160 54742 349212 54748
rect 349172 16574 349200 54742
rect 349172 16546 349292 16574
rect 348056 9172 348108 9178
rect 348056 9114 348108 9120
rect 347780 3936 347832 3942
rect 347780 3878 347832 3884
rect 348068 480 348096 9114
rect 349264 480 349292 16546
rect 350460 480 350488 60454
rect 350552 60030 351118 60058
rect 350552 6866 350580 60030
rect 353680 57730 353708 60044
rect 353668 57724 353720 57730
rect 353668 57666 353720 57672
rect 356900 57594 356928 60044
rect 356888 57588 356940 57594
rect 356888 57530 356940 57536
rect 353208 56568 353260 56574
rect 353208 56510 353260 56516
rect 351642 10296 351698 10305
rect 351642 10231 351698 10240
rect 350540 6860 350592 6866
rect 350540 6802 350592 6808
rect 351656 480 351684 10231
rect 353220 6914 353248 56510
rect 354588 53372 354640 53378
rect 354588 53314 354640 53320
rect 352852 6886 353248 6914
rect 352852 480 352880 6886
rect 354600 3398 354628 53314
rect 355232 13252 355284 13258
rect 355232 13194 355284 13200
rect 354036 3392 354088 3398
rect 354036 3334 354088 3340
rect 354588 3392 354640 3398
rect 354588 3334 354640 3340
rect 354048 480 354076 3334
rect 355244 480 355272 13194
rect 356336 5500 356388 5506
rect 356336 5442 356388 5448
rect 356348 480 356376 5442
rect 358636 5024 358688 5030
rect 358636 4966 358688 4972
rect 357532 3392 357584 3398
rect 357532 3334 357584 3340
rect 357544 480 357572 3334
rect 358648 2530 358676 4966
rect 358740 3398 358768 60454
rect 358924 60030 359490 60058
rect 361592 60030 362066 60058
rect 364444 60030 364642 60058
rect 358820 59764 358872 59770
rect 358820 59706 358872 59712
rect 358832 6914 358860 59706
rect 358924 7138 358952 60030
rect 361120 14748 361172 14754
rect 361120 14690 361172 14696
rect 358912 7132 358964 7138
rect 358912 7074 358964 7080
rect 358832 6886 359964 6914
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358648 2502 358768 2530
rect 358740 480 358768 2502
rect 359936 480 359964 6886
rect 360198 2952 360254 2961
rect 360198 2887 360200 2896
rect 360252 2887 360254 2896
rect 360200 2858 360252 2864
rect 361132 480 361160 14690
rect 361592 3738 361620 60030
rect 362868 57928 362920 57934
rect 362868 57870 362920 57876
rect 361580 3732 361632 3738
rect 361580 3674 361632 3680
rect 362880 3398 362908 57870
rect 364340 57588 364392 57594
rect 364340 57530 364392 57536
rect 363510 13152 363566 13161
rect 363510 13087 363566 13096
rect 362316 3392 362368 3398
rect 362316 3334 362368 3340
rect 362868 3392 362920 3398
rect 362868 3334 362920 3340
rect 362328 480 362356 3334
rect 363524 480 363552 13087
rect 364352 3482 364380 57530
rect 364444 4486 364472 60030
rect 367848 57594 367876 60044
rect 370424 59022 370452 60044
rect 372724 60030 373014 60058
rect 370412 59016 370464 59022
rect 370412 58958 370464 58964
rect 372620 58880 372672 58886
rect 372620 58822 372672 58828
rect 367836 57588 367888 57594
rect 367836 57530 367888 57536
rect 371148 54800 371200 54806
rect 371148 54742 371200 54748
rect 365720 53304 365772 53310
rect 365720 53246 365772 53252
rect 369768 53304 369820 53310
rect 369768 53246 369820 53252
rect 365732 16574 365760 53246
rect 367100 52080 367152 52086
rect 367100 52022 367152 52028
rect 367112 16574 367140 52022
rect 365732 16546 365852 16574
rect 367112 16546 368244 16574
rect 364432 4480 364484 4486
rect 364432 4422 364484 4428
rect 364352 3454 364656 3482
rect 364628 480 364656 3454
rect 365824 480 365852 16546
rect 367008 13184 367060 13190
rect 367008 13126 367060 13132
rect 367020 480 367048 13126
rect 368216 480 368244 16546
rect 369780 6914 369808 53246
rect 369412 6886 369808 6914
rect 369412 480 369440 6886
rect 371160 3398 371188 54742
rect 371698 9072 371754 9081
rect 371698 9007 371754 9016
rect 370596 3392 370648 3398
rect 370596 3334 370648 3340
rect 371148 3392 371200 3398
rect 371148 3334 371200 3340
rect 370608 480 370636 3334
rect 371712 480 371740 9007
rect 372632 3482 372660 58822
rect 372724 4282 372752 60030
rect 375380 59764 375432 59770
rect 375380 59706 375432 59712
rect 375288 59696 375340 59702
rect 375288 59638 375340 59644
rect 373998 10432 374054 10441
rect 373998 10367 374054 10376
rect 372712 4276 372764 4282
rect 372712 4218 372764 4224
rect 372632 3454 372936 3482
rect 372908 480 372936 3454
rect 374012 3262 374040 10367
rect 375300 3398 375328 59638
rect 375392 16574 375420 59706
rect 376220 57730 376248 60044
rect 378810 60030 379468 60058
rect 378048 59764 378100 59770
rect 378048 59706 378100 59712
rect 376208 57724 376260 57730
rect 376208 57666 376260 57672
rect 375392 16546 376524 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374000 3256 374052 3262
rect 374000 3198 374052 3204
rect 374104 480 374132 3334
rect 375288 3256 375340 3262
rect 375288 3198 375340 3204
rect 375300 480 375328 3198
rect 376496 480 376524 16546
rect 378060 6914 378088 59706
rect 378876 9036 378928 9042
rect 378876 8978 378928 8984
rect 377692 6886 378088 6914
rect 376758 2952 376814 2961
rect 376758 2887 376814 2896
rect 376772 2854 376800 2887
rect 376760 2848 376812 2854
rect 376760 2790 376812 2796
rect 377692 480 377720 6886
rect 378888 480 378916 8978
rect 379440 4486 379468 60030
rect 381372 57905 381400 60044
rect 383672 60030 383962 60058
rect 381358 57896 381414 57905
rect 381358 57831 381414 57840
rect 381544 57724 381596 57730
rect 381544 57666 381596 57672
rect 380898 18592 380954 18601
rect 380898 18527 380954 18536
rect 380912 16574 380940 18527
rect 380912 16546 381216 16574
rect 379980 14544 380032 14550
rect 379980 14486 380032 14492
rect 379428 4480 379480 4486
rect 379428 4422 379480 4428
rect 379992 480 380020 14486
rect 381188 480 381216 16546
rect 381556 13190 381584 57666
rect 382280 51876 382332 51882
rect 382280 51818 382332 51824
rect 381544 13184 381596 13190
rect 381544 13126 381596 13132
rect 382292 3398 382320 51818
rect 382372 15972 382424 15978
rect 382372 15914 382424 15920
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 15914
rect 383672 8498 383700 60030
rect 387168 57730 387196 60044
rect 387156 57724 387208 57730
rect 387156 57666 387208 57672
rect 389744 57662 389772 60044
rect 391952 60030 392334 60058
rect 394712 60030 394910 60058
rect 397472 60030 398130 60058
rect 389732 57656 389784 57662
rect 389732 57598 389784 57604
rect 386420 53236 386472 53242
rect 386420 53178 386472 53184
rect 385038 21312 385094 21321
rect 385038 21247 385094 21256
rect 385052 16574 385080 21247
rect 386432 16574 386460 53178
rect 385052 16546 386000 16574
rect 386432 16546 387196 16574
rect 384764 15904 384816 15910
rect 384764 15846 384816 15852
rect 383660 8492 383712 8498
rect 383660 8434 383712 8440
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 384776 480 384804 15846
rect 385972 480 386000 16546
rect 387168 480 387196 16546
rect 389456 14680 389508 14686
rect 389456 14622 389508 14628
rect 388260 7064 388312 7070
rect 388260 7006 388312 7012
rect 388272 480 388300 7006
rect 389468 480 389496 14622
rect 390650 11792 390706 11801
rect 390650 11727 390706 11736
rect 390664 480 390692 11727
rect 391848 7268 391900 7274
rect 391848 7210 391900 7216
rect 391860 480 391888 7210
rect 391952 5166 391980 60030
rect 393228 57180 393280 57186
rect 393228 57122 393280 57128
rect 393240 6914 393268 57122
rect 393056 6886 393268 6914
rect 391940 5160 391992 5166
rect 391940 5102 391992 5108
rect 393056 480 393084 6886
rect 394240 5160 394292 5166
rect 394240 5102 394292 5108
rect 393502 4040 393558 4049
rect 393502 3975 393558 3984
rect 393516 2990 393544 3975
rect 393504 2984 393556 2990
rect 393504 2926 393556 2932
rect 394252 480 394280 5102
rect 394712 3534 394740 60030
rect 397368 55820 397420 55826
rect 397368 55762 397420 55768
rect 395344 7336 395396 7342
rect 395344 7278 395396 7284
rect 394700 3528 394752 3534
rect 394700 3470 394752 3476
rect 395356 480 395384 7278
rect 397380 3534 397408 55762
rect 396540 3528 396592 3534
rect 396540 3470 396592 3476
rect 397368 3528 397420 3534
rect 397368 3470 397420 3476
rect 396552 480 396580 3470
rect 397472 3466 397500 60030
rect 400128 59764 400180 59770
rect 400128 59706 400180 59712
rect 400036 54936 400088 54942
rect 400036 54878 400088 54884
rect 400048 11914 400076 54878
rect 399864 11886 400076 11914
rect 399864 11694 399892 11886
rect 400140 11778 400168 59706
rect 400692 57050 400720 60044
rect 402888 58880 402940 58886
rect 402888 58822 402940 58828
rect 400680 57044 400732 57050
rect 400680 56986 400732 56992
rect 399956 11750 400168 11778
rect 399852 11688 399904 11694
rect 399852 11630 399904 11636
rect 397736 4412 397788 4418
rect 397736 4354 397788 4360
rect 397460 3460 397512 3466
rect 397460 3402 397512 3408
rect 397748 480 397776 4354
rect 399956 3534 399984 11750
rect 400128 11688 400180 11694
rect 400128 11630 400180 11636
rect 398932 3528 398984 3534
rect 398932 3470 398984 3476
rect 399944 3528 399996 3534
rect 399944 3470 399996 3476
rect 398944 480 398972 3470
rect 400140 480 400168 11630
rect 401324 10668 401376 10674
rect 401324 10610 401376 10616
rect 401336 480 401364 10610
rect 402900 6914 402928 58822
rect 403268 57662 403296 60044
rect 404268 59764 404320 59770
rect 404268 59706 404320 59712
rect 403256 57656 403308 57662
rect 403256 57598 403308 57604
rect 402532 6886 402928 6914
rect 402532 480 402560 6886
rect 404280 3534 404308 59706
rect 406488 57254 406516 60044
rect 407764 57656 407816 57662
rect 407764 57598 407816 57604
rect 406476 57248 406528 57254
rect 406476 57190 406528 57196
rect 407028 57112 407080 57118
rect 407028 57054 407080 57060
rect 407040 3534 407068 57054
rect 407212 16040 407264 16046
rect 407212 15982 407264 15988
rect 403624 3528 403676 3534
rect 403624 3470 403676 3476
rect 404268 3528 404320 3534
rect 404268 3470 404320 3476
rect 406016 3528 406068 3534
rect 406016 3470 406068 3476
rect 407028 3528 407080 3534
rect 407028 3470 407080 3476
rect 403636 480 403664 3470
rect 404820 3460 404872 3466
rect 404820 3402 404872 3408
rect 404832 480 404860 3402
rect 406028 480 406056 3470
rect 407224 480 407252 15982
rect 407776 4214 407804 57598
rect 409064 56982 409092 60044
rect 411640 57866 411668 60044
rect 414020 59696 414072 59702
rect 414020 59638 414072 59644
rect 411628 57860 411680 57866
rect 411628 57802 411680 57808
rect 409052 56976 409104 56982
rect 409052 56918 409104 56924
rect 409880 53168 409932 53174
rect 409880 53110 409932 53116
rect 409892 16574 409920 53110
rect 414032 16574 414060 59638
rect 414216 57254 414244 60044
rect 416884 60030 417450 60058
rect 414204 57248 414256 57254
rect 414204 57190 414256 57196
rect 416780 57044 416832 57050
rect 416780 56986 416832 56992
rect 409892 16546 410840 16574
rect 414032 16546 414336 16574
rect 407764 4208 407816 4214
rect 407764 4150 407816 4156
rect 409604 4208 409656 4214
rect 409604 4150 409656 4156
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 408420 480 408448 3470
rect 409616 480 409644 4150
rect 410812 480 410840 16546
rect 411904 10600 411956 10606
rect 411904 10542 411956 10548
rect 411916 480 411944 10542
rect 413100 4480 413152 4486
rect 413100 4422 413152 4428
rect 413112 480 413140 4422
rect 414308 480 414336 16546
rect 415400 14476 415452 14482
rect 415400 14418 415452 14424
rect 415412 3398 415440 14418
rect 415492 3732 415544 3738
rect 415492 3674 415544 3680
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 3674
rect 416792 3482 416820 56986
rect 416884 6526 416912 60030
rect 419540 57860 419592 57866
rect 419540 57802 419592 57808
rect 419552 16574 419580 57802
rect 420012 57050 420040 60044
rect 422404 60030 422602 60058
rect 425072 60030 425178 60058
rect 427832 60030 428398 60058
rect 430592 60030 430974 60058
rect 420920 59764 420972 59770
rect 420920 59706 420972 59712
rect 420000 57044 420052 57050
rect 420000 56986 420052 56992
rect 420932 16574 420960 59706
rect 422300 58404 422352 58410
rect 422300 58346 422352 58352
rect 419552 16546 420224 16574
rect 420932 16546 421420 16574
rect 416872 6520 416924 6526
rect 416872 6462 416924 6468
rect 418988 3936 419040 3942
rect 418988 3878 419040 3884
rect 416792 3454 417924 3482
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 417896 480 417924 3454
rect 419000 480 419028 3878
rect 420196 480 420224 16546
rect 421392 480 421420 16546
rect 422312 3482 422340 58346
rect 422404 5506 422432 60030
rect 423680 56296 423732 56302
rect 423680 56238 423732 56244
rect 423692 6914 423720 56238
rect 423772 51740 423824 51746
rect 423772 51682 423824 51688
rect 423784 11694 423812 51682
rect 423772 11688 423824 11694
rect 423772 11630 423824 11636
rect 424968 11688 425020 11694
rect 424968 11630 425020 11636
rect 423692 6886 423812 6914
rect 422392 5500 422444 5506
rect 422392 5442 422444 5448
rect 422312 3454 422616 3482
rect 422588 480 422616 3454
rect 423784 480 423812 6886
rect 424980 480 425008 11630
rect 425072 5098 425100 60030
rect 427832 6662 427860 60030
rect 429200 57044 429252 57050
rect 429200 56986 429252 56992
rect 429108 55752 429160 55758
rect 429108 55694 429160 55700
rect 427820 6656 427872 6662
rect 427820 6598 427872 6604
rect 427268 6520 427320 6526
rect 427268 6462 427320 6468
rect 425060 5092 425112 5098
rect 425060 5034 425112 5040
rect 426164 5092 426216 5098
rect 426164 5034 426216 5040
rect 426176 480 426204 5034
rect 427280 480 427308 6462
rect 429120 3398 429148 55694
rect 429212 16574 429240 56986
rect 429212 16546 429700 16574
rect 428464 3392 428516 3398
rect 428464 3334 428516 3340
rect 429108 3392 429160 3398
rect 429108 3334 429160 3340
rect 428476 480 428504 3334
rect 429672 480 429700 16546
rect 430592 5234 430620 60030
rect 431868 59628 431920 59634
rect 431868 59570 431920 59576
rect 430580 5228 430632 5234
rect 430580 5170 430632 5176
rect 431880 3398 431908 59570
rect 433536 57934 433564 60044
rect 436112 60030 436770 60058
rect 434720 58336 434772 58342
rect 434720 58278 434772 58284
rect 433524 57928 433576 57934
rect 433524 57870 433576 57876
rect 433248 56296 433300 56302
rect 433248 56238 433300 56244
rect 431960 10532 432012 10538
rect 431960 10474 432012 10480
rect 430856 3392 430908 3398
rect 430856 3334 430908 3340
rect 431868 3392 431920 3398
rect 431868 3334 431920 3340
rect 430868 480 430896 3334
rect 431972 3262 432000 10474
rect 433260 3398 433288 56238
rect 434732 16574 434760 58278
rect 436112 20670 436140 60030
rect 439332 59226 439360 60044
rect 439320 59220 439372 59226
rect 439320 59162 439372 59168
rect 439424 58478 439452 73086
rect 439502 73063 439558 73072
rect 439504 73024 439556 73030
rect 439504 72966 439556 72972
rect 439412 58472 439464 58478
rect 439412 58414 439464 58420
rect 439044 57792 439096 57798
rect 439044 57734 439096 57740
rect 436100 20664 436152 20670
rect 436100 20606 436152 20612
rect 439056 16574 439084 57734
rect 434732 16546 435588 16574
rect 439056 16546 439176 16574
rect 434444 8084 434496 8090
rect 434444 8026 434496 8032
rect 432052 3392 432104 3398
rect 432052 3334 432104 3340
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 431960 3256 432012 3262
rect 431960 3198 432012 3204
rect 432064 480 432092 3334
rect 433248 3256 433300 3262
rect 433248 3198 433300 3204
rect 433260 480 433288 3198
rect 434456 480 434484 8026
rect 435560 480 435588 16546
rect 437940 8016 437992 8022
rect 437940 7958 437992 7964
rect 436744 3324 436796 3330
rect 436744 3266 436796 3272
rect 436756 480 436784 3266
rect 437952 480 437980 7958
rect 439148 480 439176 16546
rect 439516 4554 439544 72966
rect 439608 59702 439636 152254
rect 439884 142154 439912 171106
rect 439962 166288 440018 166297
rect 439962 166223 440018 166232
rect 439700 142126 439912 142154
rect 439700 61062 439728 142126
rect 439870 96656 439926 96665
rect 439870 96591 439926 96600
rect 439778 93936 439834 93945
rect 439778 93871 439834 93880
rect 439688 61056 439740 61062
rect 439688 60998 439740 61004
rect 439596 59696 439648 59702
rect 439596 59638 439648 59644
rect 439792 53446 439820 93871
rect 439780 53440 439832 53446
rect 439780 53382 439832 53388
rect 439884 15910 439912 96591
rect 439976 54738 440004 166223
rect 440054 67688 440110 67697
rect 440054 67623 440110 67632
rect 440068 56098 440096 67623
rect 440146 64832 440202 64841
rect 440146 64767 440202 64776
rect 440056 56092 440108 56098
rect 440056 56034 440108 56040
rect 439964 54732 440016 54738
rect 439964 54674 440016 54680
rect 439872 15904 439924 15910
rect 439872 15846 439924 15852
rect 440160 5166 440188 64767
rect 440148 5160 440200 5166
rect 440148 5102 440200 5108
rect 439504 4548 439556 4554
rect 439504 4490 439556 4496
rect 440252 3398 440280 539446
rect 440344 535401 440372 656882
rect 440330 535392 440386 535401
rect 440330 535327 440386 535336
rect 440330 526552 440386 526561
rect 440330 526487 440386 526496
rect 440344 9450 440372 526487
rect 440436 521121 440464 700538
rect 447784 700460 447836 700466
rect 447784 700402 447836 700408
rect 440608 700324 440660 700330
rect 440608 700266 440660 700272
rect 442356 700324 442408 700330
rect 442356 700266 442408 700272
rect 440516 543380 440568 543386
rect 440516 543322 440568 543328
rect 440422 521112 440478 521121
rect 440422 521047 440478 521056
rect 440422 491872 440478 491881
rect 440422 491807 440478 491816
rect 440332 9444 440384 9450
rect 440332 9386 440384 9392
rect 440436 8294 440464 491807
rect 440528 61130 440556 543322
rect 440620 283121 440648 700266
rect 440792 683188 440844 683194
rect 440792 683130 440844 683136
rect 440698 451072 440754 451081
rect 440698 451007 440754 451016
rect 440606 283112 440662 283121
rect 440606 283047 440662 283056
rect 440606 242312 440662 242321
rect 440606 242247 440662 242256
rect 440516 61124 440568 61130
rect 440516 61066 440568 61072
rect 440424 8288 440476 8294
rect 440424 8230 440476 8236
rect 440620 4350 440648 242247
rect 440712 58886 440740 451007
rect 440804 427961 440832 683130
rect 442264 670744 442316 670750
rect 442264 670686 442316 670692
rect 440976 539436 441028 539442
rect 440976 539378 441028 539384
rect 440884 539096 440936 539102
rect 440884 539038 440936 539044
rect 440790 427952 440846 427961
rect 440790 427887 440846 427896
rect 440790 384432 440846 384441
rect 440790 384367 440846 384376
rect 440804 60926 440832 384367
rect 440896 365702 440924 539038
rect 440988 431934 441016 539378
rect 441068 539300 441120 539306
rect 441068 539242 441120 539248
rect 440976 431928 441028 431934
rect 440976 431870 441028 431876
rect 440884 365696 440936 365702
rect 440884 365638 440936 365644
rect 440882 306232 440938 306241
rect 440882 306167 440938 306176
rect 440792 60920 440844 60926
rect 440792 60862 440844 60868
rect 440700 58880 440752 58886
rect 440700 58822 440752 58828
rect 440896 9654 440924 306167
rect 440974 300112 441030 300121
rect 440974 300047 441030 300056
rect 440884 9648 440936 9654
rect 440884 9590 440936 9596
rect 440988 7546 441016 300047
rect 441080 259418 441108 539242
rect 442078 532672 442134 532681
rect 442078 532607 442134 532616
rect 442092 531350 442120 532607
rect 442080 531344 442132 531350
rect 442080 531286 442132 531292
rect 441618 529952 441674 529961
rect 441618 529887 441674 529896
rect 441068 259412 441120 259418
rect 441068 259354 441120 259360
rect 441066 224632 441122 224641
rect 441066 224567 441122 224576
rect 441080 57118 441108 224567
rect 441158 189952 441214 189961
rect 441158 189887 441214 189896
rect 441172 61334 441200 189887
rect 441250 183832 441306 183841
rect 441250 183767 441306 183776
rect 441264 61674 441292 183767
rect 441526 125760 441582 125769
rect 441526 125695 441582 125704
rect 441540 125662 441568 125695
rect 441528 125656 441580 125662
rect 441528 125598 441580 125604
rect 441526 122904 441582 122913
rect 441526 122839 441528 122848
rect 441580 122839 441582 122848
rect 441528 122810 441580 122816
rect 441526 119368 441582 119377
rect 441526 119303 441582 119312
rect 441540 118726 441568 119303
rect 441528 118720 441580 118726
rect 441528 118662 441580 118668
rect 441526 116648 441582 116657
rect 441526 116583 441582 116592
rect 441540 116006 441568 116583
rect 441528 116000 441580 116006
rect 441528 115942 441580 115948
rect 441526 114472 441582 114481
rect 441526 114407 441528 114416
rect 441580 114407 441582 114416
rect 441528 114378 441580 114384
rect 441526 111208 441582 111217
rect 441526 111143 441582 111152
rect 441540 110498 441568 111143
rect 441528 110492 441580 110498
rect 441528 110434 441580 110440
rect 441526 107808 441582 107817
rect 441526 107743 441582 107752
rect 441540 107710 441568 107743
rect 441528 107704 441580 107710
rect 441528 107646 441580 107652
rect 441526 105088 441582 105097
rect 441526 105023 441582 105032
rect 441540 104922 441568 105023
rect 441528 104916 441580 104922
rect 441528 104858 441580 104864
rect 441528 103488 441580 103494
rect 441526 103456 441528 103465
rect 441580 103456 441582 103465
rect 441526 103391 441582 103400
rect 441526 99648 441582 99657
rect 441526 99583 441582 99592
rect 441540 99414 441568 99583
rect 441528 99408 441580 99414
rect 441528 99350 441580 99356
rect 441526 91216 441582 91225
rect 441526 91151 441582 91160
rect 441540 91118 441568 91151
rect 441528 91112 441580 91118
rect 441528 91054 441580 91060
rect 441526 87408 441582 87417
rect 441526 87343 441582 87352
rect 441540 87038 441568 87343
rect 441528 87032 441580 87038
rect 441528 86974 441580 86980
rect 441342 85232 441398 85241
rect 441342 85167 441398 85176
rect 441252 61668 441304 61674
rect 441252 61610 441304 61616
rect 441160 61328 441212 61334
rect 441160 61270 441212 61276
rect 441356 59838 441384 85167
rect 441526 81968 441582 81977
rect 441526 81903 441582 81912
rect 441540 81462 441568 81903
rect 441528 81456 441580 81462
rect 441528 81398 441580 81404
rect 441528 80028 441580 80034
rect 441528 79970 441580 79976
rect 441540 79801 441568 79970
rect 441526 79792 441582 79801
rect 441526 79727 441582 79736
rect 441526 76392 441582 76401
rect 441526 76327 441528 76336
rect 441580 76327 441582 76336
rect 441528 76298 441580 76304
rect 441434 70952 441490 70961
rect 441434 70887 441490 70896
rect 441344 59832 441396 59838
rect 441344 59774 441396 59780
rect 441068 57112 441120 57118
rect 441068 57054 441120 57060
rect 441448 56506 441476 70887
rect 441526 61568 441582 61577
rect 441526 61503 441582 61512
rect 441540 60926 441568 61503
rect 441528 60920 441580 60926
rect 441528 60862 441580 60868
rect 441436 56500 441488 56506
rect 441436 56442 441488 56448
rect 440976 7540 441028 7546
rect 440976 7482 441028 7488
rect 440608 4344 440660 4350
rect 440608 4286 440660 4292
rect 441632 4078 441660 529887
rect 441802 500712 441858 500721
rect 441802 500647 441858 500656
rect 441816 489914 441844 500647
rect 441724 489886 441844 489914
rect 441620 4072 441672 4078
rect 441620 4014 441672 4020
rect 440332 4004 440384 4010
rect 440332 3946 440384 3952
rect 440240 3392 440292 3398
rect 440240 3334 440292 3340
rect 440344 480 440372 3946
rect 441724 3534 441752 489886
rect 441802 483032 441858 483041
rect 441802 482967 441858 482976
rect 441816 3670 441844 482967
rect 441894 477592 441950 477601
rect 441894 477527 441950 477536
rect 441908 3942 441936 477527
rect 441986 407552 442042 407561
rect 441986 407487 442042 407496
rect 441896 3936 441948 3942
rect 441896 3878 441948 3884
rect 441804 3664 441856 3670
rect 441804 3606 441856 3612
rect 441712 3528 441764 3534
rect 441712 3470 441764 3476
rect 442000 3466 442028 407487
rect 442078 402112 442134 402121
rect 442078 402047 442134 402056
rect 442092 3602 442120 402047
rect 442276 390561 442304 670686
rect 442368 442241 442396 700266
rect 442448 576904 442500 576910
rect 442448 576846 442500 576852
rect 442460 509561 442488 576846
rect 445852 543108 445904 543114
rect 445852 543050 445904 543056
rect 444380 542972 444432 542978
rect 444380 542914 444432 542920
rect 443000 539572 443052 539578
rect 443000 539514 443052 539520
rect 442538 523832 442594 523841
rect 442538 523767 442594 523776
rect 442552 523666 442580 523767
rect 442540 523660 442592 523666
rect 442540 523602 442592 523608
rect 442906 517712 442962 517721
rect 442906 517647 442962 517656
rect 442920 517546 442948 517647
rect 442908 517540 442960 517546
rect 442908 517482 442960 517488
rect 442906 514992 442962 515001
rect 442906 514927 442962 514936
rect 442920 514826 442948 514927
rect 442908 514820 442960 514826
rect 442908 514762 442960 514768
rect 442906 512272 442962 512281
rect 442906 512207 442908 512216
rect 442960 512207 442962 512216
rect 442908 512178 442960 512184
rect 442446 509552 442502 509561
rect 442446 509487 442502 509496
rect 442538 506152 442594 506161
rect 442538 506087 442594 506096
rect 442552 505170 442580 506087
rect 442540 505164 442592 505170
rect 442540 505106 442592 505112
rect 442814 503432 442870 503441
rect 442814 503367 442870 503376
rect 442828 502382 442856 503367
rect 442816 502376 442868 502382
rect 442816 502318 442868 502324
rect 442538 497992 442594 498001
rect 442538 497927 442594 497936
rect 442552 496874 442580 497927
rect 442540 496868 442592 496874
rect 442540 496810 442592 496816
rect 442722 486432 442778 486441
rect 442722 486367 442778 486376
rect 442736 485858 442764 486367
rect 442724 485852 442776 485858
rect 442724 485794 442776 485800
rect 442906 480312 442962 480321
rect 442906 480247 442908 480256
rect 442960 480247 442962 480256
rect 442908 480218 442960 480224
rect 442906 474192 442962 474201
rect 442906 474127 442962 474136
rect 442920 473414 442948 474127
rect 442908 473408 442960 473414
rect 442908 473350 442960 473356
rect 442906 471472 442962 471481
rect 442906 471407 442962 471416
rect 442920 470626 442948 471407
rect 442908 470620 442960 470626
rect 442908 470562 442960 470568
rect 442906 468752 442962 468761
rect 442906 468687 442908 468696
rect 442960 468687 442962 468696
rect 442908 468658 442960 468664
rect 442814 466032 442870 466041
rect 442814 465967 442870 465976
rect 442828 465118 442856 465967
rect 442816 465112 442868 465118
rect 442816 465054 442868 465060
rect 442906 462632 442962 462641
rect 442906 462567 442908 462576
rect 442960 462567 442962 462576
rect 442908 462538 442960 462544
rect 442906 459912 442962 459921
rect 442906 459847 442908 459856
rect 442960 459847 442962 459856
rect 442908 459818 442960 459824
rect 442906 457192 442962 457201
rect 442906 457127 442908 457136
rect 442960 457127 442962 457136
rect 442908 457098 442960 457104
rect 442906 454472 442962 454481
rect 442906 454407 442962 454416
rect 442920 454102 442948 454407
rect 442908 454096 442960 454102
rect 442908 454038 442960 454044
rect 442906 448352 442962 448361
rect 442906 448287 442962 448296
rect 442920 447506 442948 448287
rect 442908 447500 442960 447506
rect 442908 447442 442960 447448
rect 442354 442232 442410 442241
rect 442354 442167 442410 442176
rect 442722 436792 442778 436801
rect 442722 436727 442778 436736
rect 442736 436150 442764 436727
rect 442724 436144 442776 436150
rect 442724 436086 442776 436092
rect 442906 430672 442962 430681
rect 442906 430607 442908 430616
rect 442960 430607 442962 430616
rect 442908 430578 442960 430584
rect 442906 422512 442962 422521
rect 442906 422447 442962 422456
rect 442920 422346 442948 422447
rect 442908 422340 442960 422346
rect 442908 422282 442960 422288
rect 442538 419112 442594 419121
rect 442538 419047 442594 419056
rect 442552 418946 442580 419047
rect 442540 418940 442592 418946
rect 442540 418882 442592 418888
rect 442722 416392 442778 416401
rect 442722 416327 442778 416336
rect 442736 415682 442764 416327
rect 442724 415676 442776 415682
rect 442724 415618 442776 415624
rect 442538 410272 442594 410281
rect 442538 410207 442594 410216
rect 442552 409902 442580 410207
rect 442540 409896 442592 409902
rect 442540 409838 442592 409844
rect 442538 404832 442594 404841
rect 442538 404767 442594 404776
rect 442552 404666 442580 404767
rect 442540 404660 442592 404666
rect 442540 404602 442592 404608
rect 442906 395992 442962 396001
rect 442906 395927 442962 395936
rect 442920 395010 442948 395927
rect 442908 395004 442960 395010
rect 442908 394946 442960 394952
rect 442262 390552 442318 390561
rect 442262 390487 442318 390496
rect 442906 381712 442962 381721
rect 442906 381647 442962 381656
rect 442920 380934 442948 381647
rect 442908 380928 442960 380934
rect 442908 380870 442960 380876
rect 442906 378992 442962 379001
rect 442906 378927 442962 378936
rect 442920 378214 442948 378927
rect 442908 378208 442960 378214
rect 442908 378150 442960 378156
rect 442906 375592 442962 375601
rect 442906 375527 442962 375536
rect 442920 375426 442948 375527
rect 442908 375420 442960 375426
rect 442908 375362 442960 375368
rect 442906 372872 442962 372881
rect 442906 372807 442908 372816
rect 442960 372807 442962 372816
rect 442908 372778 442960 372784
rect 442170 370152 442226 370161
rect 442170 370087 442226 370096
rect 442184 4146 442212 370087
rect 442906 366752 442962 366761
rect 442906 366687 442962 366696
rect 442920 365770 442948 366687
rect 442908 365764 442960 365770
rect 442908 365706 442960 365712
rect 442630 361312 442686 361321
rect 442630 361247 442686 361256
rect 442644 360602 442672 361247
rect 442632 360596 442684 360602
rect 442632 360538 442684 360544
rect 442722 358592 442778 358601
rect 442722 358527 442778 358536
rect 442736 358426 442764 358527
rect 442724 358420 442776 358426
rect 442724 358362 442776 358368
rect 442906 355192 442962 355201
rect 442906 355127 442962 355136
rect 442920 354754 442948 355127
rect 442908 354748 442960 354754
rect 442908 354690 442960 354696
rect 442906 352472 442962 352481
rect 442906 352407 442908 352416
rect 442960 352407 442962 352416
rect 442908 352378 442960 352384
rect 442722 349752 442778 349761
rect 442722 349687 442778 349696
rect 442736 349178 442764 349687
rect 442724 349172 442776 349178
rect 442724 349114 442776 349120
rect 442906 343632 442962 343641
rect 442906 343567 442962 343576
rect 442920 342650 442948 343567
rect 442908 342644 442960 342650
rect 442908 342586 442960 342592
rect 442908 340944 442960 340950
rect 442906 340912 442908 340921
rect 442960 340912 442962 340921
rect 442906 340847 442962 340856
rect 442906 338192 442962 338201
rect 442906 338127 442908 338136
rect 442960 338127 442962 338136
rect 442908 338098 442960 338104
rect 442722 334792 442778 334801
rect 442722 334727 442778 334736
rect 442736 334218 442764 334727
rect 442724 334212 442776 334218
rect 442724 334154 442776 334160
rect 442906 332072 442962 332081
rect 442906 332007 442962 332016
rect 442920 331634 442948 332007
rect 442908 331628 442960 331634
rect 442908 331570 442960 331576
rect 442906 329352 442962 329361
rect 442906 329287 442962 329296
rect 442920 328506 442948 329287
rect 442908 328500 442960 328506
rect 442908 328442 442960 328448
rect 442538 326632 442594 326641
rect 442538 326567 442594 326576
rect 442552 326126 442580 326567
rect 442540 326120 442592 326126
rect 442540 326062 442592 326068
rect 442538 323232 442594 323241
rect 442538 323167 442594 323176
rect 442552 323134 442580 323167
rect 442540 323128 442592 323134
rect 442540 323070 442592 323076
rect 442906 320512 442962 320521
rect 442906 320447 442962 320456
rect 442920 320210 442948 320447
rect 442908 320204 442960 320210
rect 442908 320146 442960 320152
rect 442906 317792 442962 317801
rect 442906 317727 442962 317736
rect 442920 317558 442948 317727
rect 442908 317552 442960 317558
rect 442908 317494 442960 317500
rect 442262 315072 442318 315081
rect 442262 315007 442318 315016
rect 442172 4140 442224 4146
rect 442172 4082 442224 4088
rect 442080 3596 442132 3602
rect 442080 3538 442132 3544
rect 442276 3505 442304 315007
rect 442722 311672 442778 311681
rect 442722 311607 442778 311616
rect 442736 310826 442764 311607
rect 442724 310820 442776 310826
rect 442724 310762 442776 310768
rect 442906 308952 442962 308961
rect 442906 308887 442962 308896
rect 442920 307834 442948 308887
rect 442908 307828 442960 307834
rect 442908 307770 442960 307776
rect 442446 302832 442502 302841
rect 442446 302767 442502 302776
rect 442460 302530 442488 302767
rect 442448 302524 442500 302530
rect 442448 302466 442500 302472
rect 442908 298104 442960 298110
rect 442908 298046 442960 298052
rect 442920 297401 442948 298046
rect 442906 297392 442962 297401
rect 442906 297327 442962 297336
rect 442446 294672 442502 294681
rect 442446 294607 442448 294616
rect 442500 294607 442502 294616
rect 442448 294578 442500 294584
rect 442906 291272 442962 291281
rect 442906 291207 442908 291216
rect 442960 291207 442962 291216
rect 442908 291178 442960 291184
rect 442906 288552 442962 288561
rect 442906 288487 442908 288496
rect 442960 288487 442962 288496
rect 442908 288458 442960 288464
rect 442906 285832 442962 285841
rect 442906 285767 442908 285776
rect 442960 285767 442962 285776
rect 442908 285738 442960 285744
rect 442814 279712 442870 279721
rect 442814 279647 442870 279656
rect 442828 278798 442856 279647
rect 442816 278792 442868 278798
rect 442816 278734 442868 278740
rect 442538 276992 442594 277001
rect 442538 276927 442594 276936
rect 442552 276690 442580 276927
rect 442540 276684 442592 276690
rect 442540 276626 442592 276632
rect 442906 274272 442962 274281
rect 442906 274207 442962 274216
rect 442920 273290 442948 274207
rect 442908 273284 442960 273290
rect 442908 273226 442960 273232
rect 442906 271552 442962 271561
rect 442906 271487 442962 271496
rect 442920 270842 442948 271487
rect 442908 270836 442960 270842
rect 442908 270778 442960 270784
rect 442906 268152 442962 268161
rect 442906 268087 442962 268096
rect 442920 267782 442948 268087
rect 442908 267776 442960 267782
rect 442908 267718 442960 267724
rect 442906 265432 442962 265441
rect 442906 265367 442962 265376
rect 442920 264994 442948 265367
rect 442908 264988 442960 264994
rect 442908 264930 442960 264936
rect 442908 263220 442960 263226
rect 442908 263162 442960 263168
rect 442920 262721 442948 263162
rect 442906 262712 442962 262721
rect 442906 262647 442962 262656
rect 442906 259312 442962 259321
rect 442906 259247 442962 259256
rect 442920 258126 442948 259247
rect 442908 258120 442960 258126
rect 442908 258062 442960 258068
rect 442538 256592 442594 256601
rect 442538 256527 442540 256536
rect 442592 256527 442594 256536
rect 442540 256498 442592 256504
rect 442354 253872 442410 253881
rect 442354 253807 442410 253816
rect 442368 3806 442396 253807
rect 442908 251184 442960 251190
rect 442906 251152 442908 251161
rect 442960 251152 442962 251161
rect 442906 251087 442962 251096
rect 442722 247752 442778 247761
rect 442722 247687 442778 247696
rect 442736 247110 442764 247687
rect 442724 247104 442776 247110
rect 442724 247046 442776 247052
rect 442906 245032 442962 245041
rect 442906 244967 442962 244976
rect 442920 244322 442948 244967
rect 442908 244316 442960 244322
rect 442908 244258 442960 244264
rect 442722 239592 442778 239601
rect 442722 239527 442778 239536
rect 442736 239154 442764 239527
rect 442724 239148 442776 239154
rect 442724 239090 442776 239096
rect 442906 236192 442962 236201
rect 442906 236127 442962 236136
rect 442920 236026 442948 236127
rect 442908 236020 442960 236026
rect 442908 235962 442960 235968
rect 442906 233472 442962 233481
rect 442906 233407 442908 233416
rect 442960 233407 442962 233416
rect 442908 233378 442960 233384
rect 442906 230752 442962 230761
rect 442906 230687 442908 230696
rect 442960 230687 442962 230696
rect 442908 230658 442960 230664
rect 442906 227352 442962 227361
rect 442906 227287 442962 227296
rect 442920 226370 442948 227287
rect 442908 226364 442960 226370
rect 442908 226306 442960 226312
rect 442630 221912 442686 221921
rect 442630 221847 442686 221856
rect 442644 221066 442672 221847
rect 442632 221060 442684 221066
rect 442632 221002 442684 221008
rect 442906 219192 442962 219201
rect 442906 219127 442962 219136
rect 442920 218074 442948 219127
rect 442908 218068 442960 218074
rect 442908 218010 442960 218016
rect 442906 215792 442962 215801
rect 442906 215727 442962 215736
rect 442920 215354 442948 215727
rect 442908 215348 442960 215354
rect 442908 215290 442960 215296
rect 442722 213072 442778 213081
rect 442722 213007 442778 213016
rect 442736 212906 442764 213007
rect 442724 212900 442776 212906
rect 442724 212842 442776 212848
rect 442722 210352 442778 210361
rect 442722 210287 442724 210296
rect 442776 210287 442778 210296
rect 442724 210258 442776 210264
rect 442446 207632 442502 207641
rect 442446 207567 442502 207576
rect 442356 3800 442408 3806
rect 442356 3742 442408 3748
rect 442262 3496 442318 3505
rect 441988 3460 442040 3466
rect 442262 3431 442318 3440
rect 441988 3402 442040 3408
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 441540 480 441568 3334
rect 442460 3330 442488 207567
rect 442908 204264 442960 204270
rect 442906 204232 442908 204241
rect 442960 204232 442962 204241
rect 442906 204167 442962 204176
rect 442908 201544 442960 201550
rect 442906 201512 442908 201521
rect 442960 201512 442962 201521
rect 442906 201447 442962 201456
rect 442906 198792 442962 198801
rect 442906 198727 442908 198736
rect 442960 198727 442962 198736
rect 442908 198698 442960 198704
rect 442906 195392 442962 195401
rect 442906 195327 442908 195336
rect 442960 195327 442962 195336
rect 442908 195298 442960 195304
rect 442906 192672 442962 192681
rect 442906 192607 442908 192616
rect 442960 192607 442962 192616
rect 442908 192578 442960 192584
rect 442630 187232 442686 187241
rect 442630 187167 442686 187176
rect 442644 186522 442672 187167
rect 442632 186516 442684 186522
rect 442632 186458 442684 186464
rect 442906 181112 442962 181121
rect 442906 181047 442908 181056
rect 442960 181047 442962 181056
rect 442908 181018 442960 181024
rect 442906 178392 442962 178401
rect 442906 178327 442908 178336
rect 442960 178327 442962 178336
rect 442908 178298 442960 178304
rect 442722 175672 442778 175681
rect 442722 175607 442724 175616
rect 442776 175607 442778 175616
rect 442724 175578 442776 175584
rect 442906 172272 442962 172281
rect 442906 172207 442962 172216
rect 442920 171154 442948 172207
rect 442908 171148 442960 171154
rect 442908 171090 442960 171096
rect 442906 169552 442962 169561
rect 442906 169487 442962 169496
rect 442920 168434 442948 169487
rect 442908 168428 442960 168434
rect 442908 168370 442960 168376
rect 442538 164112 442594 164121
rect 442538 164047 442594 164056
rect 442552 3913 442580 164047
rect 442906 160712 442962 160721
rect 442906 160647 442908 160656
rect 442960 160647 442962 160656
rect 442908 160618 442960 160624
rect 442724 158704 442776 158710
rect 442724 158646 442776 158652
rect 442736 158001 442764 158646
rect 442722 157992 442778 158001
rect 442722 157927 442778 157936
rect 442630 155272 442686 155281
rect 442630 155207 442686 155216
rect 442538 3904 442594 3913
rect 442538 3839 442594 3848
rect 442644 3738 442672 155207
rect 442906 149152 442962 149161
rect 442906 149087 442908 149096
rect 442960 149087 442962 149096
rect 442908 149058 442960 149064
rect 442816 147620 442868 147626
rect 442816 147562 442868 147568
rect 442828 146441 442856 147562
rect 442814 146432 442870 146441
rect 442814 146367 442870 146376
rect 442906 143712 442962 143721
rect 442906 143647 442908 143656
rect 442960 143647 442962 143656
rect 442908 143618 442960 143624
rect 442906 140312 442962 140321
rect 442906 140247 442962 140256
rect 442920 139466 442948 140247
rect 442908 139460 442960 139466
rect 442908 139402 442960 139408
rect 442722 137592 442778 137601
rect 442722 137527 442778 137536
rect 442736 3777 442764 137527
rect 442906 134872 442962 134881
rect 442906 134807 442962 134816
rect 442920 132494 442948 134807
rect 442828 132466 442948 132494
rect 442722 3768 442778 3777
rect 442632 3732 442684 3738
rect 442722 3703 442778 3712
rect 442632 3674 442684 3680
rect 442632 3392 442684 3398
rect 442828 3369 442856 132466
rect 442906 132152 442962 132161
rect 442906 132087 442908 132096
rect 442960 132087 442962 132096
rect 442908 132058 442960 132064
rect 442906 128752 442962 128761
rect 442906 128687 442962 128696
rect 442920 3641 442948 128687
rect 443012 59906 443040 539514
rect 443182 413672 443238 413681
rect 443182 413607 443238 413616
rect 443090 364032 443146 364041
rect 443090 363967 443146 363976
rect 443000 59900 443052 59906
rect 443000 59842 443052 59848
rect 443104 5438 443132 363967
rect 443196 60790 443224 413607
rect 443644 360596 443696 360602
rect 443644 360538 443696 360544
rect 443552 323128 443604 323134
rect 443552 323070 443604 323076
rect 443276 302524 443328 302530
rect 443276 302466 443328 302472
rect 443184 60784 443236 60790
rect 443184 60726 443236 60732
rect 443092 5432 443144 5438
rect 443092 5374 443144 5380
rect 443288 4690 443316 302466
rect 443368 294636 443420 294642
rect 443368 294578 443420 294584
rect 443276 4684 443328 4690
rect 443276 4626 443328 4632
rect 443380 4554 443408 294578
rect 443460 276684 443512 276690
rect 443460 276626 443512 276632
rect 443472 8226 443500 276626
rect 443564 61810 443592 323070
rect 443656 245614 443684 360538
rect 443644 245608 443696 245614
rect 443644 245550 443696 245556
rect 443828 239148 443880 239154
rect 443828 239090 443880 239096
rect 443644 221060 443696 221066
rect 443644 221002 443696 221008
rect 443552 61804 443604 61810
rect 443552 61746 443604 61752
rect 443656 8566 443684 221002
rect 443736 186516 443788 186522
rect 443736 186458 443788 186464
rect 443644 8560 443696 8566
rect 443644 8502 443696 8508
rect 443460 8220 443512 8226
rect 443460 8162 443512 8168
rect 443368 4548 443420 4554
rect 443368 4490 443420 4496
rect 443748 4418 443776 186458
rect 443840 60450 443868 239090
rect 444012 212900 444064 212906
rect 444012 212842 444064 212848
rect 443920 88052 443972 88058
rect 443920 87994 443972 88000
rect 443828 60444 443880 60450
rect 443828 60386 443880 60392
rect 443932 6914 443960 87994
rect 444024 61742 444052 212842
rect 444104 114436 444156 114442
rect 444104 114378 444156 114384
rect 444012 61736 444064 61742
rect 444012 61678 444064 61684
rect 444116 61198 444144 114378
rect 444104 61192 444156 61198
rect 444104 61134 444156 61140
rect 444392 57866 444420 542914
rect 444564 352436 444616 352442
rect 444564 352378 444616 352384
rect 444472 310820 444524 310826
rect 444472 310762 444524 310768
rect 444380 57860 444432 57866
rect 444380 57802 444432 57808
rect 443840 6886 443960 6914
rect 443736 4412 443788 4418
rect 443736 4354 443788 4360
rect 442906 3632 442962 3641
rect 442906 3567 442962 3576
rect 442632 3334 442684 3340
rect 442814 3360 442870 3369
rect 442448 3324 442500 3330
rect 442448 3266 442500 3272
rect 442644 480 442672 3334
rect 442814 3295 442870 3304
rect 443840 480 443868 6886
rect 444484 6050 444512 310762
rect 444576 60586 444604 352378
rect 444656 338156 444708 338162
rect 444656 338098 444708 338104
rect 444668 60994 444696 338098
rect 445760 233436 445812 233442
rect 445760 233378 445812 233384
rect 444748 195356 444800 195362
rect 444748 195298 444800 195304
rect 444656 60988 444708 60994
rect 444656 60930 444708 60936
rect 444564 60580 444616 60586
rect 444564 60522 444616 60528
rect 444760 54942 444788 195298
rect 444840 175636 444892 175642
rect 444840 175578 444892 175584
rect 444852 60858 444880 175578
rect 444932 160676 444984 160682
rect 444932 160618 444984 160624
rect 444840 60852 444892 60858
rect 444840 60794 444892 60800
rect 444944 60518 444972 160618
rect 445024 118720 445076 118726
rect 445024 118662 445076 118668
rect 445036 88058 445064 118662
rect 445024 88052 445076 88058
rect 445024 87994 445076 88000
rect 445024 81456 445076 81462
rect 445024 81398 445076 81404
rect 444932 60512 444984 60518
rect 444932 60454 444984 60460
rect 444748 54936 444800 54942
rect 444748 54878 444800 54884
rect 445036 53582 445064 81398
rect 445116 76356 445168 76362
rect 445116 76298 445168 76304
rect 445128 55826 445156 76298
rect 445116 55820 445168 55826
rect 445116 55762 445168 55768
rect 445024 53576 445076 53582
rect 445024 53518 445076 53524
rect 445772 11762 445800 233378
rect 445864 52018 445892 543050
rect 446036 539776 446088 539782
rect 446036 539718 446088 539724
rect 445944 512236 445996 512242
rect 445944 512178 445996 512184
rect 445956 60654 445984 512178
rect 446048 103494 446076 539718
rect 447140 505164 447192 505170
rect 447140 505106 447192 505112
rect 446128 404660 446180 404666
rect 446128 404602 446180 404608
rect 446036 103488 446088 103494
rect 446036 103430 446088 103436
rect 445944 60648 445996 60654
rect 445944 60590 445996 60596
rect 446140 58954 446168 404602
rect 446312 342644 446364 342650
rect 446312 342586 446364 342592
rect 446220 334212 446272 334218
rect 446220 334154 446272 334160
rect 446128 58948 446180 58954
rect 446128 58890 446180 58896
rect 445852 52012 445904 52018
rect 445852 51954 445904 51960
rect 446128 13184 446180 13190
rect 446128 13126 446180 13132
rect 445760 11756 445812 11762
rect 445760 11698 445812 11704
rect 446140 6914 446168 13126
rect 446232 12034 446260 334154
rect 446324 61266 446352 342586
rect 446404 285796 446456 285802
rect 446404 285738 446456 285744
rect 446312 61260 446364 61266
rect 446312 61202 446364 61208
rect 446416 59974 446444 285738
rect 446496 181076 446548 181082
rect 446496 181018 446548 181024
rect 446404 59968 446456 59974
rect 446404 59910 446456 59916
rect 446508 58614 446536 181018
rect 446588 132116 446640 132122
rect 446588 132058 446640 132064
rect 446496 58608 446548 58614
rect 446496 58550 446548 58556
rect 446600 53514 446628 132058
rect 446772 122868 446824 122874
rect 446772 122810 446824 122816
rect 446680 99408 446732 99414
rect 446680 99350 446732 99356
rect 446692 55758 446720 99350
rect 446680 55752 446732 55758
rect 446680 55694 446732 55700
rect 446588 53508 446640 53514
rect 446588 53450 446640 53456
rect 446784 49026 446812 122810
rect 446772 49020 446824 49026
rect 446772 48962 446824 48968
rect 446220 12028 446272 12034
rect 446220 11970 446272 11976
rect 446140 6886 446260 6914
rect 444472 6044 444524 6050
rect 444472 5986 444524 5992
rect 445024 4208 445076 4214
rect 445024 4150 445076 4156
rect 445036 480 445064 4150
rect 446232 480 446260 6886
rect 447152 5370 447180 505106
rect 447508 496868 447560 496874
rect 447508 496810 447560 496816
rect 447232 462596 447284 462602
rect 447232 462538 447284 462544
rect 447244 6118 447272 462538
rect 447416 459876 447468 459882
rect 447416 459818 447468 459824
rect 447324 457156 447376 457162
rect 447324 457098 447376 457104
rect 447232 6112 447284 6118
rect 447232 6054 447284 6060
rect 447336 5982 447364 457098
rect 447428 8634 447456 459818
rect 447520 50454 447548 496810
rect 447600 468716 447652 468722
rect 447600 468658 447652 468664
rect 447612 56234 447640 468658
rect 447692 415676 447744 415682
rect 447692 415618 447744 415624
rect 447600 56228 447652 56234
rect 447600 56170 447652 56176
rect 447508 50448 447560 50454
rect 447508 50390 447560 50396
rect 447416 8628 447468 8634
rect 447416 8570 447468 8576
rect 447324 5976 447376 5982
rect 447324 5918 447376 5924
rect 447140 5364 447192 5370
rect 447140 5306 447192 5312
rect 447704 5098 447732 415618
rect 447796 263226 447824 700402
rect 449900 697604 449952 697610
rect 449900 697546 449952 697552
rect 448612 543176 448664 543182
rect 448612 543118 448664 543124
rect 448520 523660 448572 523666
rect 448520 523602 448572 523608
rect 447876 358420 447928 358426
rect 447876 358362 447928 358368
rect 447784 263220 447836 263226
rect 447784 263162 447836 263168
rect 447784 57316 447836 57322
rect 447784 57258 447836 57264
rect 447692 5092 447744 5098
rect 447692 5034 447744 5040
rect 447796 3482 447824 57258
rect 447888 8702 447916 358362
rect 447968 331628 448020 331634
rect 447968 331570 448020 331576
rect 447980 60382 448008 331570
rect 448060 291236 448112 291242
rect 448060 291178 448112 291184
rect 447968 60376 448020 60382
rect 447968 60318 448020 60324
rect 448072 58818 448100 291178
rect 448244 270836 448296 270842
rect 448244 270778 448296 270784
rect 448152 256556 448204 256562
rect 448152 256498 448204 256504
rect 448164 60246 448192 256498
rect 448256 60314 448284 270778
rect 448244 60308 448296 60314
rect 448244 60250 448296 60256
rect 448152 60240 448204 60246
rect 448152 60182 448204 60188
rect 448060 58812 448112 58818
rect 448060 58754 448112 58760
rect 447876 8696 447928 8702
rect 447876 8638 447928 8644
rect 448532 6390 448560 523602
rect 448624 59770 448652 543118
rect 448704 447500 448756 447506
rect 448704 447442 448756 447448
rect 448612 59764 448664 59770
rect 448612 59706 448664 59712
rect 448612 57248 448664 57254
rect 448612 57190 448664 57196
rect 448520 6384 448572 6390
rect 448520 6326 448572 6332
rect 448520 4820 448572 4826
rect 448520 4762 448572 4768
rect 447428 3454 447824 3482
rect 447428 480 447456 3454
rect 448532 2394 448560 4762
rect 448624 3534 448652 57190
rect 448716 10742 448744 447442
rect 448796 430636 448848 430642
rect 448796 430578 448848 430584
rect 448808 39438 448836 430578
rect 448888 395004 448940 395010
rect 448888 394946 448940 394952
rect 448796 39432 448848 39438
rect 448796 39374 448848 39380
rect 448704 10736 448756 10742
rect 448704 10678 448756 10684
rect 448900 6730 448928 394946
rect 448980 372836 449032 372842
rect 448980 372778 449032 372784
rect 448888 6724 448940 6730
rect 448888 6666 448940 6672
rect 448992 6458 449020 372778
rect 449072 317552 449124 317558
rect 449072 317494 449124 317500
rect 449084 60178 449112 317494
rect 449164 230716 449216 230722
rect 449164 230658 449216 230664
rect 449072 60172 449124 60178
rect 449072 60114 449124 60120
rect 448980 6452 449032 6458
rect 448980 6394 449032 6400
rect 449176 6322 449204 230658
rect 449256 143676 449308 143682
rect 449256 143618 449308 143624
rect 449268 57186 449296 143618
rect 449912 80034 449940 697546
rect 450084 543312 450136 543318
rect 450084 543254 450136 543260
rect 449992 542904 450044 542910
rect 449992 542846 450044 542852
rect 449900 80028 449952 80034
rect 449900 79970 449952 79976
rect 449256 57180 449308 57186
rect 449256 57122 449308 57128
rect 449900 10464 449952 10470
rect 449900 10406 449952 10412
rect 449164 6316 449216 6322
rect 449164 6258 449216 6264
rect 448612 3528 448664 3534
rect 448612 3470 448664 3476
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 449912 3482 449940 10406
rect 450004 4214 450032 542846
rect 450096 58410 450124 543254
rect 452660 542836 452712 542842
rect 452660 542778 452712 542784
rect 451280 514820 451332 514826
rect 451280 514762 451332 514768
rect 450176 418940 450228 418946
rect 450176 418882 450228 418888
rect 450084 58404 450136 58410
rect 450084 58346 450136 58352
rect 450188 14618 450216 418882
rect 450268 326120 450320 326126
rect 450268 326062 450320 326068
rect 450176 14612 450228 14618
rect 450176 14554 450228 14560
rect 450280 11830 450308 326062
rect 450360 288516 450412 288522
rect 450360 288458 450412 288464
rect 450372 11898 450400 288458
rect 450452 210316 450504 210322
rect 450452 210258 450504 210264
rect 450464 56370 450492 210258
rect 450544 192636 450596 192642
rect 450544 192578 450596 192584
rect 450452 56364 450504 56370
rect 450452 56306 450504 56312
rect 450556 53310 450584 192578
rect 450636 178356 450688 178362
rect 450636 178298 450688 178304
rect 450648 56438 450676 178298
rect 451292 56574 451320 514762
rect 451372 320204 451424 320210
rect 451372 320146 451424 320152
rect 451280 56568 451332 56574
rect 451280 56510 451332 56516
rect 450636 56432 450688 56438
rect 450636 56374 450688 56380
rect 451384 54874 451412 320146
rect 451556 244316 451608 244322
rect 451556 244258 451608 244264
rect 451464 110492 451516 110498
rect 451464 110434 451516 110440
rect 451372 54868 451424 54874
rect 451372 54810 451424 54816
rect 450544 53304 450596 53310
rect 450544 53246 450596 53252
rect 451476 16574 451504 110434
rect 451568 55078 451596 244258
rect 451648 168428 451700 168434
rect 451648 168370 451700 168376
rect 451556 55072 451608 55078
rect 451556 55014 451608 55020
rect 451660 51950 451688 168370
rect 452672 58342 452700 542778
rect 454132 542700 454184 542706
rect 454132 542642 454184 542648
rect 454040 541272 454092 541278
rect 454040 541214 454092 541220
rect 452752 470620 452804 470626
rect 452752 470562 452804 470568
rect 452660 58336 452712 58342
rect 452660 58278 452712 58284
rect 451648 51944 451700 51950
rect 451648 51886 451700 51892
rect 451476 16546 452148 16574
rect 450360 11892 450412 11898
rect 450360 11834 450412 11840
rect 450268 11824 450320 11830
rect 450268 11766 450320 11772
rect 449992 4208 450044 4214
rect 449992 4150 450044 4156
rect 448532 2366 448652 2394
rect 448624 480 448652 2366
rect 449820 480 449848 3470
rect 449912 3454 450952 3482
rect 450924 480 450952 3454
rect 452120 480 452148 16546
rect 452764 11966 452792 470562
rect 452844 454096 452896 454102
rect 452844 454038 452896 454044
rect 452856 13326 452884 454038
rect 452936 422340 452988 422346
rect 452936 422282 452988 422288
rect 452948 54806 452976 422282
rect 453028 236020 453080 236026
rect 453028 235962 453080 235968
rect 452936 54800 452988 54806
rect 452936 54742 452988 54748
rect 453040 26926 453068 235962
rect 453120 198756 453172 198762
rect 453120 198698 453172 198704
rect 453132 53378 453160 198698
rect 453120 53372 453172 53378
rect 453120 53314 453172 53320
rect 453028 26920 453080 26926
rect 453028 26862 453080 26868
rect 452844 13320 452896 13326
rect 452844 13262 452896 13268
rect 452752 11960 452804 11966
rect 452752 11902 452804 11908
rect 454052 3398 454080 541214
rect 454144 6526 454172 542642
rect 456984 541612 457036 541618
rect 456984 541554 457036 541560
rect 456800 541000 456852 541006
rect 456800 540942 456852 540948
rect 455420 539912 455472 539918
rect 455420 539854 455472 539860
rect 454684 480276 454736 480282
rect 454684 480218 454736 480224
rect 454224 328500 454276 328506
rect 454224 328442 454276 328448
rect 454236 56302 454264 328442
rect 454316 267776 454368 267782
rect 454316 267718 454368 267724
rect 454224 56296 454276 56302
rect 454224 56238 454276 56244
rect 454328 22846 454356 267718
rect 454408 247104 454460 247110
rect 454408 247046 454460 247052
rect 454420 50522 454448 247046
rect 454696 113150 454724 480218
rect 454684 113144 454736 113150
rect 454684 113086 454736 113092
rect 454408 50516 454460 50522
rect 454408 50458 454460 50464
rect 454316 22840 454368 22846
rect 454316 22782 454368 22788
rect 454132 6520 454184 6526
rect 454132 6462 454184 6468
rect 455432 4010 455460 539854
rect 455696 5296 455748 5302
rect 455696 5238 455748 5244
rect 455420 4004 455472 4010
rect 455420 3946 455472 3952
rect 454500 3868 454552 3874
rect 454500 3810 454552 3816
rect 454040 3392 454092 3398
rect 454040 3334 454092 3340
rect 453304 3188 453356 3194
rect 453304 3130 453356 3136
rect 453316 480 453344 3130
rect 454512 480 454540 3810
rect 455708 480 455736 5238
rect 456812 3482 456840 540942
rect 456892 473408 456944 473414
rect 456892 473350 456944 473356
rect 456904 3602 456932 473350
rect 456892 3596 456944 3602
rect 456892 3538 456944 3544
rect 456812 3454 456932 3482
rect 456904 480 456932 3454
rect 456996 3194 457024 541554
rect 458824 541136 458876 541142
rect 458824 541078 458876 541084
rect 457076 409896 457128 409902
rect 457076 409838 457128 409844
rect 457088 50590 457116 409838
rect 457076 50584 457128 50590
rect 457076 50526 457128 50532
rect 458088 3596 458140 3602
rect 458088 3538 458140 3544
rect 456984 3188 457036 3194
rect 456984 3130 457036 3136
rect 458100 480 458128 3538
rect 458836 3534 458864 541078
rect 461584 340944 461636 340950
rect 461584 340886 461636 340892
rect 460204 139460 460256 139466
rect 460204 139402 460256 139408
rect 459192 7472 459244 7478
rect 459192 7414 459244 7420
rect 458824 3528 458876 3534
rect 458824 3470 458876 3476
rect 459204 480 459232 7414
rect 460216 4554 460244 139402
rect 461596 6914 461624 340886
rect 461676 91112 461728 91118
rect 461676 91054 461728 91060
rect 461504 6886 461624 6914
rect 460204 4548 460256 4554
rect 460204 4490 460256 4496
rect 460388 3528 460440 3534
rect 460388 3470 460440 3476
rect 460400 480 460428 3470
rect 461504 3466 461532 6886
rect 461688 6866 461716 91054
rect 462332 58546 462360 703520
rect 478524 700534 478552 703520
rect 464344 700528 464396 700534
rect 464344 700470 464396 700476
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 464356 204270 464384 700470
rect 494808 698970 494836 703520
rect 527192 700466 527220 703520
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543476 700330 543504 703520
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 494796 698964 494848 698970
rect 494796 698906 494848 698912
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579618 591016 579674 591025
rect 579618 590951 579674 590960
rect 579632 590714 579660 590951
rect 579620 590708 579672 590714
rect 579620 590650 579672 590656
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 475384 543040 475436 543046
rect 475384 542982 475436 542988
rect 468484 540116 468536 540122
rect 468484 540058 468536 540064
rect 466460 537940 466512 537946
rect 466460 537882 466512 537888
rect 465724 307828 465776 307834
rect 465724 307770 465776 307776
rect 464344 204264 464396 204270
rect 464344 204206 464396 204212
rect 465080 125656 465132 125662
rect 465080 125598 465132 125604
rect 462320 58540 462372 58546
rect 462320 58482 462372 58488
rect 463700 57724 463752 57730
rect 463700 57666 463752 57672
rect 463712 16574 463740 57666
rect 465092 16574 465120 125598
rect 463712 16546 464016 16574
rect 465092 16546 465212 16574
rect 461676 6860 461728 6866
rect 461676 6802 461728 6808
rect 461584 6792 461636 6798
rect 461584 6734 461636 6740
rect 461492 3460 461544 3466
rect 461492 3402 461544 3408
rect 461596 480 461624 6734
rect 462780 4548 462832 4554
rect 462780 4490 462832 4496
rect 462792 480 462820 4490
rect 463988 480 464016 16546
rect 465184 480 465212 16546
rect 465736 3534 465764 307770
rect 466472 16574 466500 537882
rect 466472 16546 467512 16574
rect 466276 7880 466328 7886
rect 466276 7822 466328 7828
rect 465724 3528 465776 3534
rect 465724 3470 465776 3476
rect 466288 480 466316 7822
rect 467484 480 467512 16546
rect 468392 10396 468444 10402
rect 468392 10338 468444 10344
rect 468404 3482 468432 10338
rect 468496 3670 468524 540058
rect 472624 258120 472676 258126
rect 472624 258062 472676 258068
rect 470600 53100 470652 53106
rect 470600 53042 470652 53048
rect 470612 16574 470640 53042
rect 472636 33114 472664 258062
rect 472716 56160 472768 56166
rect 472716 56102 472768 56108
rect 472624 33108 472676 33114
rect 472624 33050 472676 33056
rect 470612 16546 471100 16574
rect 469864 7812 469916 7818
rect 469864 7754 469916 7760
rect 468484 3664 468536 3670
rect 468484 3606 468536 3612
rect 468404 3454 468708 3482
rect 468680 480 468708 3454
rect 469876 480 469904 7754
rect 471072 480 471100 16546
rect 472728 3534 472756 56102
rect 475396 4554 475424 542982
rect 511264 542768 511316 542774
rect 511264 542710 511316 542716
rect 498844 542632 498896 542638
rect 498844 542574 498896 542580
rect 479524 541544 479576 541550
rect 479524 541486 479576 541492
rect 477500 104916 477552 104922
rect 477500 104858 477552 104864
rect 476120 39364 476172 39370
rect 476120 39306 476172 39312
rect 476132 16574 476160 39306
rect 477512 16574 477540 104858
rect 476132 16546 476988 16574
rect 477512 16546 478184 16574
rect 475384 4548 475436 4554
rect 475384 4490 475436 4496
rect 474556 3664 474608 3670
rect 474556 3606 474608 3612
rect 473452 3596 473504 3602
rect 473452 3538 473504 3544
rect 472716 3528 472768 3534
rect 472716 3470 472768 3476
rect 472254 3224 472310 3233
rect 472254 3159 472310 3168
rect 472268 480 472296 3159
rect 473464 480 473492 3538
rect 474568 480 474596 3606
rect 475752 3528 475804 3534
rect 475752 3470 475804 3476
rect 475764 480 475792 3470
rect 476960 480 476988 16546
rect 478156 480 478184 16546
rect 479340 10328 479392 10334
rect 479340 10270 479392 10276
rect 479352 480 479380 10270
rect 479536 3534 479564 541486
rect 486424 541408 486476 541414
rect 486424 541350 486476 541356
rect 483020 538824 483072 538830
rect 483020 538766 483072 538772
rect 481640 531344 481692 531350
rect 481640 531286 481692 531292
rect 480260 226364 480312 226370
rect 480260 226306 480312 226312
rect 480272 16574 480300 226306
rect 480272 16546 480576 16574
rect 479524 3528 479576 3534
rect 479524 3470 479576 3476
rect 480548 480 480576 16546
rect 481652 3602 481680 531286
rect 483032 16574 483060 538766
rect 485044 264988 485096 264994
rect 485044 264930 485096 264936
rect 484400 61600 484452 61606
rect 484400 61542 484452 61548
rect 484412 16574 484440 61542
rect 483032 16546 484072 16574
rect 484412 16546 484992 16574
rect 481732 4548 481784 4554
rect 481732 4490 481784 4496
rect 481640 3596 481692 3602
rect 481640 3538 481692 3544
rect 481744 480 481772 4490
rect 482836 3596 482888 3602
rect 482836 3538 482888 3544
rect 482848 480 482876 3538
rect 484044 480 484072 16546
rect 484964 3482 484992 16546
rect 485056 4078 485084 264930
rect 485780 50380 485832 50386
rect 485780 50322 485832 50328
rect 485792 6914 485820 50322
rect 486436 16574 486464 541350
rect 493324 540048 493376 540054
rect 493324 539990 493376 539996
rect 487160 538348 487212 538354
rect 487160 538290 487212 538296
rect 487172 16574 487200 538290
rect 490012 502376 490064 502382
rect 490012 502318 490064 502324
rect 488540 61532 488592 61538
rect 488540 61474 488592 61480
rect 488552 16574 488580 61474
rect 490024 16574 490052 502318
rect 492680 47592 492732 47598
rect 492680 47534 492732 47540
rect 492692 16574 492720 47534
rect 486436 16546 486556 16574
rect 487172 16546 487660 16574
rect 488552 16546 488856 16574
rect 490024 16546 491156 16574
rect 492692 16546 493272 16574
rect 485792 6886 486464 6914
rect 485044 4072 485096 4078
rect 485044 4014 485096 4020
rect 484964 3454 485268 3482
rect 485240 480 485268 3454
rect 486436 480 486464 6886
rect 486528 3602 486556 16546
rect 486516 3596 486568 3602
rect 486516 3538 486568 3544
rect 487632 480 487660 16546
rect 488828 480 488856 16546
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 489932 480 489960 3470
rect 491128 480 491156 16546
rect 492312 4072 492364 4078
rect 492312 4014 492364 4020
rect 492324 480 492352 4014
rect 493244 3482 493272 16546
rect 493336 3806 493364 539990
rect 498200 378208 498252 378214
rect 498200 378150 498252 378156
rect 496820 354748 496872 354754
rect 496820 354690 496872 354696
rect 494704 116000 494756 116006
rect 494704 115942 494756 115948
rect 494716 16574 494744 115942
rect 496832 16574 496860 354690
rect 494716 16546 494836 16574
rect 496832 16546 497136 16574
rect 494704 13116 494756 13122
rect 494704 13058 494756 13064
rect 493324 3800 493376 3806
rect 493324 3742 493376 3748
rect 493244 3454 493548 3482
rect 493520 480 493548 3454
rect 494716 480 494744 13058
rect 494808 3738 494836 16546
rect 494796 3732 494848 3738
rect 494796 3674 494848 3680
rect 495900 3460 495952 3466
rect 495900 3402 495952 3408
rect 495912 480 495940 3402
rect 497108 480 497136 16546
rect 498212 480 498240 378150
rect 498292 61464 498344 61470
rect 498292 61406 498344 61412
rect 498304 16574 498332 61406
rect 498304 16546 498792 16574
rect 498764 3482 498792 16546
rect 498856 3670 498884 542574
rect 503720 542496 503772 542502
rect 503720 542438 503772 542444
rect 499580 541068 499632 541074
rect 499580 541010 499632 541016
rect 499592 16574 499620 541010
rect 502340 539708 502392 539714
rect 502340 539650 502392 539656
rect 500960 149116 501012 149122
rect 500960 149058 501012 149064
rect 500224 17264 500276 17270
rect 500224 17206 500276 17212
rect 499592 16546 500172 16574
rect 498844 3664 498896 3670
rect 498844 3606 498896 3612
rect 500144 3482 500172 16546
rect 500236 3874 500264 17206
rect 500972 16574 501000 149058
rect 502352 16574 502380 539650
rect 503732 16574 503760 542438
rect 505100 538960 505152 538966
rect 505100 538902 505152 538908
rect 505112 16574 505140 538902
rect 508504 375420 508556 375426
rect 508504 375362 508556 375368
rect 506572 349172 506624 349178
rect 506572 349114 506624 349120
rect 506584 16574 506612 349114
rect 508516 219434 508544 375362
rect 508504 219428 508556 219434
rect 508504 219370 508556 219376
rect 507860 218068 507912 218074
rect 507860 218010 507912 218016
rect 507124 60920 507176 60926
rect 507124 60862 507176 60868
rect 500972 16546 501828 16574
rect 502352 16546 503024 16574
rect 503732 16546 504220 16574
rect 505112 16546 505416 16574
rect 506584 16546 507072 16574
rect 500224 3868 500276 3874
rect 500224 3810 500276 3816
rect 498764 3454 499436 3482
rect 500144 3454 500632 3482
rect 499408 480 499436 3454
rect 500604 480 500632 3454
rect 501800 480 501828 16546
rect 502996 480 503024 16546
rect 504192 480 504220 16546
rect 505388 480 505416 16546
rect 506480 3868 506532 3874
rect 506480 3810 506532 3816
rect 506492 480 506520 3810
rect 507044 3346 507072 16546
rect 507136 3466 507164 60862
rect 507872 16574 507900 218010
rect 509240 61396 509292 61402
rect 509240 61338 509292 61344
rect 509252 16574 509280 61338
rect 509884 57452 509936 57458
rect 509884 57394 509936 57400
rect 507872 16546 508912 16574
rect 509252 16546 509832 16574
rect 507124 3460 507176 3466
rect 507124 3402 507176 3408
rect 507044 3318 507716 3346
rect 507688 480 507716 3318
rect 508884 480 508912 16546
rect 509804 3346 509832 16546
rect 509896 3534 509924 57394
rect 511276 4826 511304 542710
rect 522304 541476 522356 541482
rect 522304 541418 522356 541424
rect 518164 541204 518216 541210
rect 518164 541146 518216 541152
rect 513380 539980 513432 539986
rect 513380 539922 513432 539928
rect 512000 539232 512052 539238
rect 512000 539174 512052 539180
rect 512012 16574 512040 539174
rect 513392 16574 513420 539922
rect 516784 436144 516836 436150
rect 516784 436086 516836 436092
rect 515404 107704 515456 107710
rect 515404 107646 515456 107652
rect 512012 16546 512500 16574
rect 513392 16546 513604 16574
rect 511264 4820 511316 4826
rect 511264 4762 511316 4768
rect 511264 3800 511316 3806
rect 511264 3742 511316 3748
rect 509884 3528 509936 3534
rect 509884 3470 509936 3476
rect 509804 3318 510108 3346
rect 510080 480 510108 3318
rect 511276 480 511304 3742
rect 512472 480 512500 16546
rect 513576 480 513604 16546
rect 515416 10334 515444 107646
rect 515404 10328 515456 10334
rect 515404 10270 515456 10276
rect 515956 6248 516008 6254
rect 515956 6190 516008 6196
rect 514760 3596 514812 3602
rect 514760 3538 514812 3544
rect 514772 480 514800 3538
rect 515968 480 515996 6190
rect 516796 3534 516824 436086
rect 517152 7948 517204 7954
rect 517152 7890 517204 7896
rect 516784 3528 516836 3534
rect 516784 3470 516836 3476
rect 517164 480 517192 7890
rect 518176 3874 518204 541146
rect 518900 380928 518952 380934
rect 518900 380870 518952 380876
rect 518256 57588 518308 57594
rect 518256 57530 518308 57536
rect 518164 3868 518216 3874
rect 518164 3810 518216 3816
rect 518268 3806 518296 57530
rect 518912 16574 518940 380870
rect 520924 278792 520976 278798
rect 520924 278734 520976 278740
rect 518912 16546 519584 16574
rect 518256 3800 518308 3806
rect 518256 3742 518308 3748
rect 518348 3528 518400 3534
rect 518348 3470 518400 3476
rect 518360 480 518388 3470
rect 519556 480 519584 16546
rect 520740 4820 520792 4826
rect 520740 4762 520792 4768
rect 520752 480 520780 4762
rect 520936 4010 520964 278734
rect 520924 4004 520976 4010
rect 520924 3946 520976 3952
rect 521844 3800 521896 3806
rect 521844 3742 521896 3748
rect 521856 480 521884 3742
rect 522316 3602 522344 541418
rect 566464 541340 566516 541346
rect 566464 541282 566516 541288
rect 531412 539844 531464 539850
rect 531412 539786 531464 539792
rect 529940 539164 529992 539170
rect 529940 539106 529992 539112
rect 527824 517540 527876 517546
rect 527824 517482 527876 517488
rect 525800 171148 525852 171154
rect 525800 171090 525852 171096
rect 524420 58744 524472 58750
rect 524420 58686 524472 58692
rect 523684 57384 523736 57390
rect 523684 57326 523736 57332
rect 523040 6180 523092 6186
rect 523040 6122 523092 6128
rect 522304 3596 522356 3602
rect 522304 3538 522356 3544
rect 523052 480 523080 6122
rect 523696 3942 523724 57326
rect 524432 16574 524460 58686
rect 525812 16574 525840 171090
rect 527180 56024 527232 56030
rect 527180 55966 527232 55972
rect 524432 16546 525472 16574
rect 525812 16546 526668 16574
rect 523684 3936 523736 3942
rect 523684 3878 523736 3884
rect 524236 3596 524288 3602
rect 524236 3538 524288 3544
rect 524248 480 524276 3538
rect 525444 480 525472 16546
rect 526640 480 526668 16546
rect 527192 6914 527220 55966
rect 527836 16574 527864 517482
rect 529204 273284 529256 273290
rect 529204 273226 529256 273232
rect 528560 25560 528612 25566
rect 528560 25502 528612 25508
rect 528572 16574 528600 25502
rect 527836 16546 527956 16574
rect 528572 16546 529060 16574
rect 527192 6886 527864 6914
rect 527836 480 527864 6886
rect 527928 3806 527956 16546
rect 527916 3800 527968 3806
rect 527916 3742 527968 3748
rect 529032 480 529060 16546
rect 529216 4078 529244 273226
rect 529952 16574 529980 539106
rect 529952 16546 530164 16574
rect 529204 4072 529256 4078
rect 529204 4014 529256 4020
rect 530136 480 530164 16546
rect 531424 6914 531452 539786
rect 556252 539640 556304 539646
rect 556252 539582 556304 539588
rect 543740 539368 543792 539374
rect 543740 539310 543792 539316
rect 539692 538484 539744 538490
rect 539692 538426 539744 538432
rect 533344 485852 533396 485858
rect 533344 485794 533396 485800
rect 531964 57520 532016 57526
rect 531964 57462 532016 57468
rect 531332 6886 531452 6914
rect 531332 480 531360 6886
rect 531976 4010 532004 57462
rect 533356 4214 533384 485794
rect 538864 465112 538916 465118
rect 538864 465054 538916 465060
rect 537484 201544 537536 201550
rect 537484 201486 537536 201492
rect 536104 28280 536156 28286
rect 536104 28222 536156 28228
rect 533712 4888 533764 4894
rect 533712 4830 533764 4836
rect 533344 4208 533396 4214
rect 533344 4150 533396 4156
rect 531964 4004 532016 4010
rect 531964 3946 532016 3952
rect 532516 3868 532568 3874
rect 532516 3810 532568 3816
rect 532528 480 532556 3810
rect 533724 480 533752 4830
rect 534908 4208 534960 4214
rect 534908 4150 534960 4156
rect 534920 480 534948 4150
rect 536116 4146 536144 28222
rect 537208 4956 537260 4962
rect 537208 4898 537260 4904
rect 536104 4140 536156 4146
rect 536104 4082 536156 4088
rect 536104 3936 536156 3942
rect 536104 3878 536156 3884
rect 536116 480 536144 3878
rect 537220 480 537248 4898
rect 537496 4894 537524 201486
rect 537484 4888 537536 4894
rect 537484 4830 537536 4836
rect 538404 4888 538456 4894
rect 538404 4830 538456 4836
rect 538416 480 538444 4830
rect 538876 3942 538904 465054
rect 539704 16574 539732 538426
rect 543004 57656 543056 57662
rect 543004 57598 543056 57604
rect 540980 54664 541032 54670
rect 540980 54606 541032 54612
rect 540992 16574 541020 54606
rect 539704 16546 540836 16574
rect 540992 16546 542032 16574
rect 539600 4140 539652 4146
rect 539600 4082 539652 4088
rect 538864 3936 538916 3942
rect 538864 3878 538916 3884
rect 539612 480 539640 4082
rect 540808 480 540836 16546
rect 542004 480 542032 16546
rect 543016 3874 543044 57598
rect 543752 16574 543780 539310
rect 550640 539028 550692 539034
rect 550640 538970 550692 538976
rect 547880 365764 547932 365770
rect 547880 365706 547932 365712
rect 545764 215348 545816 215354
rect 545764 215290 545816 215296
rect 543752 16546 544424 16574
rect 543004 3868 543056 3874
rect 543004 3810 543056 3816
rect 543188 3800 543240 3806
rect 543188 3742 543240 3748
rect 543200 480 543228 3742
rect 544396 480 544424 16546
rect 545488 8152 545540 8158
rect 545488 8094 545540 8100
rect 545500 480 545528 8094
rect 545776 3806 545804 215290
rect 546684 4072 546736 4078
rect 546684 4014 546736 4020
rect 545764 3800 545816 3806
rect 545764 3742 545816 3748
rect 546696 480 546724 4014
rect 547892 480 547920 365706
rect 548524 87032 548576 87038
rect 548524 86974 548576 86980
rect 548536 2922 548564 86974
rect 549260 60104 549312 60110
rect 549260 60046 549312 60052
rect 549272 16574 549300 60046
rect 550652 16574 550680 538970
rect 555424 51808 555476 51814
rect 555424 51750 555476 51756
rect 549272 16546 550312 16574
rect 550652 16546 551508 16574
rect 549076 7744 549128 7750
rect 549076 7686 549128 7692
rect 548524 2916 548576 2922
rect 548524 2858 548576 2864
rect 549088 480 549116 7686
rect 550284 480 550312 16546
rect 551480 480 551508 16546
rect 553768 4004 553820 4010
rect 553768 3946 553820 3952
rect 552664 3732 552716 3738
rect 552664 3674 552716 3680
rect 552676 480 552704 3674
rect 553780 480 553808 3946
rect 555436 3398 555464 51750
rect 556264 6914 556292 539582
rect 566476 100706 566504 541282
rect 580172 538892 580224 538898
rect 580172 538834 580224 538840
rect 580080 538416 580132 538422
rect 580080 538358 580132 538364
rect 579988 431928 580040 431934
rect 579988 431870 580040 431876
rect 580000 431633 580028 431870
rect 579986 431624 580042 431633
rect 579986 431559 580042 431568
rect 579988 365696 580040 365702
rect 579988 365638 580040 365644
rect 580000 365129 580028 365638
rect 579986 365120 580042 365129
rect 579986 365055 580042 365064
rect 580092 351937 580120 538358
rect 580078 351928 580134 351937
rect 580078 351863 580134 351872
rect 580184 325281 580212 538834
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 219428 580040 219434
rect 579988 219370 580040 219376
rect 580000 219065 580028 219370
rect 579986 219056 580042 219065
rect 579986 218991 580042 219000
rect 579988 113144 580040 113150
rect 579988 113086 580040 113092
rect 580000 112849 580028 113086
rect 579986 112840 580042 112849
rect 579986 112775 580042 112784
rect 566464 100700 566516 100706
rect 566464 100642 566516 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 560298 61432 560354 61441
rect 560298 61367 560354 61376
rect 557540 54596 557592 54602
rect 557540 54538 557592 54544
rect 557552 16574 557580 54538
rect 560312 16574 560340 61367
rect 567200 60036 567252 60042
rect 567200 59978 567252 59984
rect 564532 58676 564584 58682
rect 564532 58618 564584 58624
rect 564544 16574 564572 58618
rect 567212 16574 567240 59978
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580184 59430 580212 59599
rect 580172 59424 580224 59430
rect 580172 59366 580224 59372
rect 580276 59294 580304 683839
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580264 59288 580316 59294
rect 580264 59230 580316 59236
rect 580368 59022 580396 643991
rect 580540 538756 580592 538762
rect 580540 538698 580592 538704
rect 580448 538280 580500 538286
rect 580448 538222 580500 538228
rect 580460 471481 580488 538222
rect 580446 471472 580502 471481
rect 580446 471407 580502 471416
rect 580446 458144 580502 458153
rect 580446 458079 580502 458088
rect 580460 59362 580488 458079
rect 580552 152697 580580 538698
rect 580908 538688 580960 538694
rect 580908 538630 580960 538636
rect 580724 538620 580776 538626
rect 580724 538562 580776 538568
rect 580632 538552 580684 538558
rect 580632 538494 580684 538500
rect 580644 165889 580672 538494
rect 580736 537849 580764 538562
rect 580920 538214 580948 538630
rect 580828 538186 580948 538214
rect 580722 537840 580778 537849
rect 580722 537775 580778 537784
rect 580828 533338 580856 538186
rect 580908 537804 580960 537810
rect 580908 537746 580960 537752
rect 580736 533310 580856 533338
rect 580736 272241 580764 533310
rect 580920 528554 580948 537746
rect 580828 528526 580948 528554
rect 580828 524521 580856 528526
rect 580814 524512 580870 524521
rect 580814 524447 580870 524456
rect 580906 511320 580962 511329
rect 580906 511255 580962 511264
rect 580814 484664 580870 484673
rect 580814 484599 580870 484608
rect 580722 272232 580778 272241
rect 580722 272167 580778 272176
rect 580828 251190 580856 484599
rect 580920 298110 580948 511255
rect 580908 298104 580960 298110
rect 580908 298046 580960 298052
rect 580816 251184 580868 251190
rect 580816 251126 580868 251132
rect 580814 205728 580870 205737
rect 580814 205663 580870 205672
rect 580722 192536 580778 192545
rect 580722 192471 580778 192480
rect 580630 165880 580686 165889
rect 580630 165815 580686 165824
rect 580538 152688 580594 152697
rect 580538 152623 580594 152632
rect 580538 86184 580594 86193
rect 580538 86119 580594 86128
rect 580552 60722 580580 86119
rect 580736 74534 580764 192471
rect 580828 158710 580856 205663
rect 580906 179208 580962 179217
rect 580906 179143 580962 179152
rect 580816 158704 580868 158710
rect 580816 158646 580868 158652
rect 580920 147626 580948 179143
rect 580908 147620 580960 147626
rect 580908 147562 580960 147568
rect 580736 74506 580856 74534
rect 580630 72992 580686 73001
rect 580630 72927 580686 72936
rect 580540 60716 580592 60722
rect 580540 60658 580592 60664
rect 580448 59356 580500 59362
rect 580448 59298 580500 59304
rect 580644 59158 580672 72927
rect 580632 59152 580684 59158
rect 580632 59094 580684 59100
rect 580828 59090 580856 74506
rect 580816 59084 580868 59090
rect 580816 59026 580868 59032
rect 580356 59016 580408 59022
rect 580356 58958 580408 58964
rect 568580 55956 568632 55962
rect 568580 55898 568632 55904
rect 568592 16574 568620 55898
rect 580264 55888 580316 55894
rect 580264 55830 580316 55836
rect 575480 54528 575532 54534
rect 575480 54470 575532 54476
rect 575492 16574 575520 54470
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580276 19825 580304 55830
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 557552 16546 558592 16574
rect 560312 16546 560892 16574
rect 564544 16546 565676 16574
rect 567212 16546 568068 16574
rect 568592 16546 569172 16574
rect 575492 16546 576348 16574
rect 556172 6886 556292 6914
rect 555424 3392 555476 3398
rect 555424 3334 555476 3340
rect 554964 2916 555016 2922
rect 554964 2858 555016 2864
rect 554976 480 555004 2858
rect 556172 480 556200 6886
rect 557356 3392 557408 3398
rect 557356 3334 557408 3340
rect 557368 480 557396 3334
rect 558564 480 558592 16546
rect 559748 3664 559800 3670
rect 559748 3606 559800 3612
rect 559760 480 559788 3606
rect 560864 480 560892 16546
rect 562048 10328 562100 10334
rect 562048 10270 562100 10276
rect 562060 480 562088 10270
rect 563242 7576 563298 7585
rect 563242 7511 563298 7520
rect 563256 480 563284 7511
rect 564440 3936 564492 3942
rect 564440 3878 564492 3884
rect 564452 480 564480 3878
rect 565648 480 565676 16546
rect 566832 7676 566884 7682
rect 566832 7618 566884 7624
rect 566844 480 566872 7618
rect 568040 480 568068 16546
rect 569144 480 569172 16546
rect 571524 8968 571576 8974
rect 571524 8910 571576 8916
rect 570328 3460 570380 3466
rect 570328 3402 570380 3408
rect 570340 480 570368 3402
rect 571536 480 571564 8910
rect 572720 5024 572772 5030
rect 572720 4966 572772 4972
rect 572732 480 572760 4966
rect 575112 3868 575164 3874
rect 575112 3810 575164 3816
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 573928 480 573956 3470
rect 575124 480 575152 3810
rect 576320 480 576348 16546
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 577424 480 577452 7550
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581000 6588 581052 6594
rect 581000 6530 581052 6536
rect 578608 3800 578660 3806
rect 578608 3742 578660 3748
rect 578620 480 578648 3742
rect 581012 480 581040 6530
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 582208 480 582236 3538
rect 583390 3088 583446 3097
rect 583390 3023 583446 3032
rect 583404 480 583432 3023
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632032 3478 632088
rect 3238 527856 3294 527912
rect 3330 514800 3386 514856
rect 3790 619112 3846 619168
rect 3606 606056 3662 606112
rect 3514 579944 3570 580000
rect 3514 566888 3570 566944
rect 3330 501744 3386 501800
rect 3422 475632 3478 475688
rect 3422 410488 3478 410544
rect 3330 319232 3386 319288
rect 2778 254108 2834 254144
rect 2778 254088 2780 254108
rect 2780 254088 2832 254108
rect 2832 254088 2834 254108
rect 3054 241032 3110 241088
rect 3146 202816 3202 202872
rect 3146 201864 3202 201920
rect 3330 188808 3386 188864
rect 2778 149776 2834 149832
rect 3330 136720 3386 136776
rect 3146 111696 3202 111752
rect 3146 110608 3202 110664
rect 3330 84632 3386 84688
rect 2962 58520 3018 58576
rect 3698 553832 3754 553888
rect 3698 423544 3754 423600
rect 3606 398656 3662 398712
rect 3606 397432 3662 397488
rect 3606 371320 3662 371376
rect 3514 214920 3570 214976
rect 3514 71576 3570 71632
rect 3698 358400 3754 358456
rect 3790 345344 3846 345400
rect 3974 449520 4030 449576
rect 3974 293120 4030 293176
rect 3882 267144 3938 267200
rect 3882 162832 3938 162888
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 32408 3478 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 23018 3304 23074 3360
rect 34794 3440 34850 3496
rect 40682 3576 40738 3632
rect 45466 3712 45522 3768
rect 53102 61376 53158 61432
rect 54758 7520 54814 7576
rect 56506 506776 56562 506832
rect 56414 442856 56470 442912
rect 56322 440136 56378 440192
rect 56230 408176 56286 408232
rect 56046 355816 56102 355872
rect 55954 335416 56010 335472
rect 55862 280336 55918 280392
rect 56138 326576 56194 326632
rect 56598 268776 56654 268832
rect 56598 216416 56654 216472
rect 56598 198756 56654 198792
rect 56598 198736 56600 198756
rect 56600 198736 56652 198756
rect 56652 198736 56654 198756
rect 56598 103556 56654 103592
rect 56598 103536 56600 103556
rect 56600 103536 56652 103556
rect 56652 103536 56654 103556
rect 57426 529932 57428 529952
rect 57428 529932 57480 529952
rect 57480 529932 57482 529952
rect 57426 529896 57482 529932
rect 57334 527196 57390 527232
rect 57334 527176 57336 527196
rect 57336 527176 57388 527196
rect 57388 527176 57390 527196
rect 57334 524476 57390 524512
rect 57334 524456 57336 524476
rect 57336 524456 57388 524476
rect 57388 524456 57390 524476
rect 57334 521056 57390 521112
rect 57334 518336 57390 518392
rect 57334 515616 57390 515672
rect 57334 512896 57390 512952
rect 57150 509496 57206 509552
rect 57058 477556 57114 477592
rect 57058 477536 57060 477556
rect 57060 477536 57112 477556
rect 57112 477536 57114 477556
rect 56874 465976 56930 466032
rect 57058 445576 57114 445632
rect 56874 367376 56930 367432
rect 56874 364656 56930 364712
rect 56874 350376 56930 350432
rect 57334 323856 57390 323912
rect 56874 315016 56930 315072
rect 57334 312296 57390 312352
rect 57334 309576 57390 309632
rect 57334 300736 57390 300792
rect 57334 298016 57390 298072
rect 57058 291896 57114 291952
rect 57334 289176 57390 289232
rect 57334 283056 57390 283112
rect 57334 277616 57390 277672
rect 57334 271496 57390 271552
rect 57518 504056 57574 504112
rect 57610 495216 57666 495272
rect 57610 492496 57666 492552
rect 57610 489096 57666 489152
rect 57610 480936 57666 480992
rect 57610 474816 57666 474872
rect 57610 469376 57666 469432
rect 57610 463256 57666 463312
rect 57610 460536 57666 460592
rect 57610 457816 57666 457872
rect 57610 454416 57666 454472
rect 57610 451696 57666 451752
rect 57610 437416 57666 437472
rect 57610 434016 57666 434072
rect 57610 431296 57666 431352
rect 57610 428576 57666 428632
rect 57610 422456 57666 422512
rect 57610 419736 57666 419792
rect 57610 417016 57666 417072
rect 57610 413616 57666 413672
rect 57518 410896 57574 410952
rect 57518 402056 57574 402112
rect 57518 399336 57574 399392
rect 57518 396616 57574 396672
rect 57518 393896 57574 393952
rect 57518 390496 57574 390552
rect 57518 387812 57520 387832
rect 57520 387812 57572 387832
rect 57572 387812 57574 387832
rect 57518 387776 57574 387812
rect 57518 385076 57574 385112
rect 57518 385056 57520 385076
rect 57520 385056 57572 385076
rect 57572 385056 57574 385076
rect 57518 381656 57574 381712
rect 57518 378936 57574 378992
rect 57518 373496 57574 373552
rect 57518 361936 57574 361992
rect 57518 358536 57574 358592
rect 57518 353096 57574 353152
rect 57518 346976 57574 347032
rect 57518 341536 57574 341592
rect 57518 338156 57574 338192
rect 57518 338136 57520 338156
rect 57520 338136 57572 338156
rect 57572 338136 57574 338156
rect 57518 329976 57574 330032
rect 57426 266056 57482 266112
rect 57426 262656 57482 262712
rect 57334 259936 57390 259992
rect 57426 254496 57482 254552
rect 56874 251096 56930 251152
rect 57426 248376 57482 248432
rect 57334 242956 57390 242992
rect 57334 242936 57336 242956
rect 57336 242936 57388 242956
rect 57388 242936 57390 242956
rect 57334 239536 57390 239592
rect 57242 234096 57298 234152
rect 56874 190576 56930 190632
rect 57150 158616 57206 158672
rect 57058 143656 57114 143712
rect 56966 126656 57022 126712
rect 56874 77016 56930 77072
rect 56782 71576 56838 71632
rect 56874 65456 56930 65512
rect 57334 230696 57390 230752
rect 57242 3032 57298 3088
rect 59082 533296 59138 533352
rect 57794 483656 57850 483712
rect 58990 472096 59046 472152
rect 57794 448976 57850 449032
rect 58898 405456 58954 405512
rect 58806 376216 58862 376272
rect 57886 332696 57942 332752
rect 57978 321136 58034 321192
rect 57886 294616 57942 294672
rect 57886 236816 57942 236872
rect 57886 227976 57942 228032
rect 57886 225256 57942 225312
rect 57886 222536 57942 222592
rect 57886 219136 57942 219192
rect 57886 210976 57942 211032
rect 57702 207576 57758 207632
rect 57702 204856 57758 204912
rect 57702 196036 57758 196072
rect 57702 196016 57704 196036
rect 57704 196016 57756 196036
rect 57756 196016 57758 196036
rect 57702 193296 57758 193352
rect 57702 187176 57758 187232
rect 57702 184456 57758 184512
rect 57702 181736 57758 181792
rect 57702 172896 57758 172952
rect 57886 202136 57942 202192
rect 57886 175616 57942 175672
rect 57886 170176 57942 170232
rect 57886 166776 57942 166832
rect 57886 164056 57942 164112
rect 57886 155216 57942 155272
rect 57886 152496 57942 152552
rect 57886 149776 57942 149832
rect 57886 147056 57942 147112
rect 57886 140936 57942 140992
rect 57886 135496 57942 135552
rect 57886 132096 57942 132152
rect 57886 129376 57942 129432
rect 57886 123256 57942 123312
rect 57886 120536 57942 120592
rect 57886 117816 57942 117872
rect 57886 115096 57942 115152
rect 57886 106256 57942 106312
rect 57886 100136 57942 100192
rect 57886 94696 57942 94752
rect 57886 88576 57942 88632
rect 57886 85856 57942 85912
rect 58714 286456 58770 286512
rect 58622 257216 58678 257272
rect 58530 245656 58586 245712
rect 58438 97416 58494 97472
rect 58346 91296 58402 91352
rect 58254 83136 58310 83192
rect 58162 74296 58218 74352
rect 58070 68176 58126 68232
rect 59174 501336 59230 501392
rect 113454 542544 113510 542600
rect 132774 543496 132830 543552
rect 218978 699760 219034 699816
rect 226798 543632 226854 543688
rect 146942 542816 146998 542872
rect 138570 542408 138626 542464
rect 149518 542544 149574 542600
rect 168838 543088 168894 543144
rect 166262 542952 166318 543008
rect 179786 543360 179842 543416
rect 177210 542408 177266 542464
rect 190734 542408 190790 542464
rect 210054 542544 210110 542600
rect 215206 541184 215262 541240
rect 231950 542408 232006 542464
rect 251270 542544 251326 542600
rect 257066 542408 257122 542464
rect 292486 543224 292542 543280
rect 347226 543088 347282 543144
rect 311806 542952 311862 543008
rect 336278 542680 336334 542736
rect 358818 542816 358874 542872
rect 353022 542544 353078 542600
rect 366546 542544 366602 542600
rect 391662 542816 391718 542872
rect 380714 542680 380770 542736
rect 396814 542544 396870 542600
rect 410982 542952 411038 543008
rect 72606 539552 72662 539608
rect 75642 539552 75698 539608
rect 106094 539552 106150 539608
rect 116306 539552 116362 539608
rect 119526 539552 119582 539608
rect 125322 539552 125378 539608
rect 127346 539552 127402 539608
rect 155590 539552 155646 539608
rect 220634 539552 220690 539608
rect 243174 539552 243230 539608
rect 253570 539552 253626 539608
rect 283838 539552 283894 539608
rect 314106 539552 314162 539608
rect 330850 539552 330906 539608
rect 341706 539552 341762 539608
rect 361026 539552 361082 539608
rect 377310 539552 377366 539608
rect 382922 539552 382978 539608
rect 385498 539552 385554 539608
rect 388810 539552 388866 539608
rect 393962 539552 394018 539608
rect 402242 539552 402298 539608
rect 60646 539436 60702 539472
rect 60646 539416 60648 539436
rect 60648 539416 60700 539436
rect 60700 539416 60702 539436
rect 223486 539416 223542 539472
rect 240230 539416 240286 539472
rect 270314 539416 270370 539472
rect 278870 539416 278926 539472
rect 298190 539416 298246 539472
rect 309138 539416 309194 539472
rect 350354 539416 350410 539472
rect 59818 536560 59874 536616
rect 59358 497936 59414 497992
rect 59266 138216 59322 138272
rect 59266 108976 59322 109032
rect 59450 425856 59506 425912
rect 59542 318416 59598 318472
rect 59634 306176 59690 306232
rect 439502 445848 439558 445904
rect 439502 438912 439558 438968
rect 439962 537920 440018 537976
rect 439870 495080 439926 495136
rect 439778 387640 439834 387696
rect 439502 152360 439558 152416
rect 59726 111696 59782 111752
rect 59818 79736 59874 79792
rect 59818 62736 59874 62792
rect 60830 2760 60886 2816
rect 64326 3848 64382 3904
rect 66718 2760 66774 2816
rect 71686 3032 71742 3088
rect 71594 2760 71650 2816
rect 73802 3168 73858 3224
rect 92754 2760 92810 2816
rect 109314 3984 109370 4040
rect 108118 3032 108174 3088
rect 106922 2896 106978 2952
rect 110510 2896 110566 2952
rect 117594 3984 117650 4040
rect 118790 3032 118846 3088
rect 137926 21256 137982 21312
rect 139306 12960 139362 13016
rect 144826 24112 144882 24168
rect 145930 11600 145986 11656
rect 155866 17448 155922 17504
rect 154210 7656 154266 7712
rect 162766 21392 162822 21448
rect 193218 4120 193274 4176
rect 205546 11736 205602 11792
rect 217966 18672 218022 18728
rect 216586 12008 216642 12064
rect 231766 14592 231822 14648
rect 237378 26832 237434 26888
rect 235814 4120 235870 4176
rect 240506 14456 240562 14512
rect 244094 5616 244150 5672
rect 246394 15816 246450 15872
rect 252466 24112 252522 24168
rect 253478 10920 253534 10976
rect 261758 5616 261814 5672
rect 281538 17312 281594 17368
rect 276018 4120 276074 4176
rect 279514 4120 279570 4176
rect 293682 10376 293738 10432
rect 296626 15816 296682 15872
rect 305550 3032 305606 3088
rect 307850 11872 307906 11928
rect 322938 17176 322994 17232
rect 332506 15816 332562 15872
rect 329838 3052 329894 3088
rect 329838 3032 329840 3052
rect 329840 3032 329892 3052
rect 329892 3032 329894 3052
rect 336278 9560 336334 9616
rect 332690 5616 332746 5672
rect 333886 4120 333942 4176
rect 342166 40568 342222 40624
rect 344558 8880 344614 8936
rect 351642 10240 351698 10296
rect 360198 2916 360254 2952
rect 360198 2896 360200 2916
rect 360200 2896 360252 2916
rect 360252 2896 360254 2916
rect 363510 13096 363566 13152
rect 371698 9016 371754 9072
rect 373998 10376 374054 10432
rect 376758 2896 376814 2952
rect 381358 57840 381414 57896
rect 380898 18536 380954 18592
rect 385038 21256 385094 21312
rect 390650 11736 390706 11792
rect 393502 3984 393558 4040
rect 439502 73072 439558 73128
rect 439962 166232 440018 166288
rect 439870 96600 439926 96656
rect 439778 93880 439834 93936
rect 440054 67632 440110 67688
rect 440146 64776 440202 64832
rect 440330 535336 440386 535392
rect 440330 526496 440386 526552
rect 440422 521056 440478 521112
rect 440422 491816 440478 491872
rect 440698 451016 440754 451072
rect 440606 283056 440662 283112
rect 440606 242256 440662 242312
rect 440790 427896 440846 427952
rect 440790 384376 440846 384432
rect 440882 306176 440938 306232
rect 440974 300056 441030 300112
rect 442078 532616 442134 532672
rect 441618 529896 441674 529952
rect 441066 224576 441122 224632
rect 441158 189896 441214 189952
rect 441250 183776 441306 183832
rect 441526 125704 441582 125760
rect 441526 122868 441582 122904
rect 441526 122848 441528 122868
rect 441528 122848 441580 122868
rect 441580 122848 441582 122868
rect 441526 119312 441582 119368
rect 441526 116592 441582 116648
rect 441526 114436 441582 114472
rect 441526 114416 441528 114436
rect 441528 114416 441580 114436
rect 441580 114416 441582 114436
rect 441526 111152 441582 111208
rect 441526 107752 441582 107808
rect 441526 105032 441582 105088
rect 441526 103436 441528 103456
rect 441528 103436 441580 103456
rect 441580 103436 441582 103456
rect 441526 103400 441582 103436
rect 441526 99592 441582 99648
rect 441526 91160 441582 91216
rect 441526 87352 441582 87408
rect 441342 85176 441398 85232
rect 441526 81912 441582 81968
rect 441526 79736 441582 79792
rect 441526 76356 441582 76392
rect 441526 76336 441528 76356
rect 441528 76336 441580 76356
rect 441580 76336 441582 76356
rect 441434 70896 441490 70952
rect 441526 61512 441582 61568
rect 441802 500656 441858 500712
rect 441802 482976 441858 483032
rect 441894 477536 441950 477592
rect 441986 407496 442042 407552
rect 442078 402056 442134 402112
rect 442538 523776 442594 523832
rect 442906 517656 442962 517712
rect 442906 514936 442962 514992
rect 442906 512236 442962 512272
rect 442906 512216 442908 512236
rect 442908 512216 442960 512236
rect 442960 512216 442962 512236
rect 442446 509496 442502 509552
rect 442538 506096 442594 506152
rect 442814 503376 442870 503432
rect 442538 497936 442594 497992
rect 442722 486376 442778 486432
rect 442906 480276 442962 480312
rect 442906 480256 442908 480276
rect 442908 480256 442960 480276
rect 442960 480256 442962 480276
rect 442906 474136 442962 474192
rect 442906 471416 442962 471472
rect 442906 468716 442962 468752
rect 442906 468696 442908 468716
rect 442908 468696 442960 468716
rect 442960 468696 442962 468716
rect 442814 465976 442870 466032
rect 442906 462596 442962 462632
rect 442906 462576 442908 462596
rect 442908 462576 442960 462596
rect 442960 462576 442962 462596
rect 442906 459876 442962 459912
rect 442906 459856 442908 459876
rect 442908 459856 442960 459876
rect 442960 459856 442962 459876
rect 442906 457156 442962 457192
rect 442906 457136 442908 457156
rect 442908 457136 442960 457156
rect 442960 457136 442962 457156
rect 442906 454416 442962 454472
rect 442906 448296 442962 448352
rect 442354 442176 442410 442232
rect 442722 436736 442778 436792
rect 442906 430636 442962 430672
rect 442906 430616 442908 430636
rect 442908 430616 442960 430636
rect 442960 430616 442962 430636
rect 442906 422456 442962 422512
rect 442538 419056 442594 419112
rect 442722 416336 442778 416392
rect 442538 410216 442594 410272
rect 442538 404776 442594 404832
rect 442906 395936 442962 395992
rect 442262 390496 442318 390552
rect 442906 381656 442962 381712
rect 442906 378936 442962 378992
rect 442906 375536 442962 375592
rect 442906 372836 442962 372872
rect 442906 372816 442908 372836
rect 442908 372816 442960 372836
rect 442960 372816 442962 372836
rect 442170 370096 442226 370152
rect 442906 366696 442962 366752
rect 442630 361256 442686 361312
rect 442722 358536 442778 358592
rect 442906 355136 442962 355192
rect 442906 352436 442962 352472
rect 442906 352416 442908 352436
rect 442908 352416 442960 352436
rect 442960 352416 442962 352436
rect 442722 349696 442778 349752
rect 442906 343576 442962 343632
rect 442906 340892 442908 340912
rect 442908 340892 442960 340912
rect 442960 340892 442962 340912
rect 442906 340856 442962 340892
rect 442906 338156 442962 338192
rect 442906 338136 442908 338156
rect 442908 338136 442960 338156
rect 442960 338136 442962 338156
rect 442722 334736 442778 334792
rect 442906 332016 442962 332072
rect 442906 329296 442962 329352
rect 442538 326576 442594 326632
rect 442538 323176 442594 323232
rect 442906 320456 442962 320512
rect 442906 317736 442962 317792
rect 442262 315016 442318 315072
rect 442722 311616 442778 311672
rect 442906 308896 442962 308952
rect 442446 302776 442502 302832
rect 442906 297336 442962 297392
rect 442446 294636 442502 294672
rect 442446 294616 442448 294636
rect 442448 294616 442500 294636
rect 442500 294616 442502 294636
rect 442906 291236 442962 291272
rect 442906 291216 442908 291236
rect 442908 291216 442960 291236
rect 442960 291216 442962 291236
rect 442906 288516 442962 288552
rect 442906 288496 442908 288516
rect 442908 288496 442960 288516
rect 442960 288496 442962 288516
rect 442906 285796 442962 285832
rect 442906 285776 442908 285796
rect 442908 285776 442960 285796
rect 442960 285776 442962 285796
rect 442814 279656 442870 279712
rect 442538 276936 442594 276992
rect 442906 274216 442962 274272
rect 442906 271496 442962 271552
rect 442906 268096 442962 268152
rect 442906 265376 442962 265432
rect 442906 262656 442962 262712
rect 442906 259256 442962 259312
rect 442538 256556 442594 256592
rect 442538 256536 442540 256556
rect 442540 256536 442592 256556
rect 442592 256536 442594 256556
rect 442354 253816 442410 253872
rect 442906 251132 442908 251152
rect 442908 251132 442960 251152
rect 442960 251132 442962 251152
rect 442906 251096 442962 251132
rect 442722 247696 442778 247752
rect 442906 244976 442962 245032
rect 442722 239536 442778 239592
rect 442906 236136 442962 236192
rect 442906 233436 442962 233472
rect 442906 233416 442908 233436
rect 442908 233416 442960 233436
rect 442960 233416 442962 233436
rect 442906 230716 442962 230752
rect 442906 230696 442908 230716
rect 442908 230696 442960 230716
rect 442960 230696 442962 230716
rect 442906 227296 442962 227352
rect 442630 221856 442686 221912
rect 442906 219136 442962 219192
rect 442906 215736 442962 215792
rect 442722 213016 442778 213072
rect 442722 210316 442778 210352
rect 442722 210296 442724 210316
rect 442724 210296 442776 210316
rect 442776 210296 442778 210316
rect 442446 207576 442502 207632
rect 442262 3440 442318 3496
rect 442906 204212 442908 204232
rect 442908 204212 442960 204232
rect 442960 204212 442962 204232
rect 442906 204176 442962 204212
rect 442906 201492 442908 201512
rect 442908 201492 442960 201512
rect 442960 201492 442962 201512
rect 442906 201456 442962 201492
rect 442906 198756 442962 198792
rect 442906 198736 442908 198756
rect 442908 198736 442960 198756
rect 442960 198736 442962 198756
rect 442906 195356 442962 195392
rect 442906 195336 442908 195356
rect 442908 195336 442960 195356
rect 442960 195336 442962 195356
rect 442906 192636 442962 192672
rect 442906 192616 442908 192636
rect 442908 192616 442960 192636
rect 442960 192616 442962 192636
rect 442630 187176 442686 187232
rect 442906 181076 442962 181112
rect 442906 181056 442908 181076
rect 442908 181056 442960 181076
rect 442960 181056 442962 181076
rect 442906 178356 442962 178392
rect 442906 178336 442908 178356
rect 442908 178336 442960 178356
rect 442960 178336 442962 178356
rect 442722 175636 442778 175672
rect 442722 175616 442724 175636
rect 442724 175616 442776 175636
rect 442776 175616 442778 175636
rect 442906 172216 442962 172272
rect 442906 169496 442962 169552
rect 442538 164056 442594 164112
rect 442906 160676 442962 160712
rect 442906 160656 442908 160676
rect 442908 160656 442960 160676
rect 442960 160656 442962 160676
rect 442722 157936 442778 157992
rect 442630 155216 442686 155272
rect 442538 3848 442594 3904
rect 442906 149116 442962 149152
rect 442906 149096 442908 149116
rect 442908 149096 442960 149116
rect 442960 149096 442962 149116
rect 442814 146376 442870 146432
rect 442906 143676 442962 143712
rect 442906 143656 442908 143676
rect 442908 143656 442960 143676
rect 442960 143656 442962 143676
rect 442906 140256 442962 140312
rect 442722 137536 442778 137592
rect 442906 134816 442962 134872
rect 442722 3712 442778 3768
rect 442906 132116 442962 132152
rect 442906 132096 442908 132116
rect 442908 132096 442960 132116
rect 442960 132096 442962 132116
rect 442906 128696 442962 128752
rect 443182 413616 443238 413672
rect 443090 363976 443146 364032
rect 442906 3576 442962 3632
rect 442814 3304 442870 3360
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579618 590960 579674 591016
rect 579618 577632 579674 577688
rect 579894 564304 579950 564360
rect 472254 3168 472310 3224
rect 579986 431568 580042 431624
rect 579986 365064 580042 365120
rect 580078 351872 580134 351928
rect 580170 325216 580226 325272
rect 579802 258848 579858 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 219000 580042 219056
rect 579986 112784 580042 112840
rect 580170 99456 580226 99512
rect 560298 61376 560354 61432
rect 580170 59608 580226 59664
rect 580354 644000 580410 644056
rect 580446 471416 580502 471472
rect 580446 458088 580502 458144
rect 580722 537784 580778 537840
rect 580814 524456 580870 524512
rect 580906 511264 580962 511320
rect 580814 484608 580870 484664
rect 580722 272176 580778 272232
rect 580814 205672 580870 205728
rect 580722 192480 580778 192536
rect 580630 165824 580686 165880
rect 580538 152632 580594 152688
rect 580538 86128 580594 86184
rect 580906 179152 580962 179208
rect 580630 72936 580686 72992
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580262 19760 580318 19816
rect 563242 7520 563298 7576
rect 580170 6568 580226 6624
rect 583390 3032 583446 3088
<< metal3 >>
rect 218973 699818 219039 699821
rect 219198 699818 219204 699820
rect 218973 699816 219204 699818
rect 218973 699760 218978 699816
rect 219034 699760 219204 699816
rect 218973 699758 219204 699760
rect 218973 699755 219039 699758
rect 219198 699756 219204 699758
rect 219268 699756 219274 699820
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3785 619170 3851 619173
rect -960 619168 3851 619170
rect -960 619112 3790 619168
rect 3846 619112 3851 619168
rect -960 619110 3851 619112
rect -960 619020 480 619110
rect 3785 619107 3851 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579613 591018 579679 591021
rect 583520 591018 584960 591108
rect 579613 591016 584960 591018
rect 579613 590960 579618 591016
rect 579674 590960 584960 591016
rect 579613 590958 584960 590960
rect 579613 590955 579679 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3693 553890 3759 553893
rect -960 553888 3759 553890
rect -960 553832 3698 553888
rect 3754 553832 3759 553888
rect -960 553830 3759 553832
rect -960 553740 480 553830
rect 3693 553827 3759 553830
rect 583520 551020 584960 551260
rect 226793 543690 226859 543693
rect 251766 543690 251772 543692
rect 226793 543688 251772 543690
rect 226793 543632 226798 543688
rect 226854 543632 251772 543688
rect 226793 543630 251772 543632
rect 226793 543627 226859 543630
rect 251766 543628 251772 543630
rect 251836 543628 251842 543692
rect 132769 543554 132835 543557
rect 277894 543554 277900 543556
rect 132769 543552 277900 543554
rect 132769 543496 132774 543552
rect 132830 543496 277900 543552
rect 132769 543494 277900 543496
rect 132769 543491 132835 543494
rect 277894 543492 277900 543494
rect 277964 543492 277970 543556
rect 179781 543418 179847 543421
rect 327574 543418 327580 543420
rect 179781 543416 327580 543418
rect 179781 543360 179786 543416
rect 179842 543360 327580 543416
rect 179781 543358 327580 543360
rect 179781 543355 179847 543358
rect 327574 543356 327580 543358
rect 327644 543356 327650 543420
rect 228214 543220 228220 543284
rect 228284 543282 228290 543284
rect 292481 543282 292547 543285
rect 228284 543280 292547 543282
rect 228284 543224 292486 543280
rect 292542 543224 292547 543280
rect 228284 543222 292547 543224
rect 228284 543220 228290 543222
rect 292481 543219 292547 543222
rect 168833 543146 168899 543149
rect 230974 543146 230980 543148
rect 168833 543144 230980 543146
rect 168833 543088 168838 543144
rect 168894 543088 230980 543144
rect 168833 543086 230980 543088
rect 168833 543083 168899 543086
rect 230974 543084 230980 543086
rect 231044 543084 231050 543148
rect 255814 543084 255820 543148
rect 255884 543146 255890 543148
rect 347221 543146 347287 543149
rect 255884 543144 347287 543146
rect 255884 543088 347226 543144
rect 347282 543088 347287 543144
rect 255884 543086 347287 543088
rect 255884 543084 255890 543086
rect 347221 543083 347287 543086
rect 166257 543010 166323 543013
rect 280654 543010 280660 543012
rect 166257 543008 280660 543010
rect 166257 542952 166262 543008
rect 166318 542952 280660 543008
rect 166257 542950 280660 542952
rect 166257 542947 166323 542950
rect 280654 542948 280660 542950
rect 280724 542948 280730 543012
rect 311801 543010 311867 543013
rect 331806 543010 331812 543012
rect 311801 543008 331812 543010
rect 311801 542952 311806 543008
rect 311862 542952 331812 543008
rect 311801 542950 331812 542952
rect 311801 542947 311867 542950
rect 331806 542948 331812 542950
rect 331876 542948 331882 543012
rect 335854 542948 335860 543012
rect 335924 543010 335930 543012
rect 410977 543010 411043 543013
rect 335924 543008 411043 543010
rect 335924 542952 410982 543008
rect 411038 542952 411043 543008
rect 335924 542950 411043 542952
rect 335924 542948 335930 542950
rect 410977 542947 411043 542950
rect 146937 542874 147003 542877
rect 271086 542874 271092 542876
rect 146937 542872 271092 542874
rect 146937 542816 146942 542872
rect 146998 542816 271092 542872
rect 146937 542814 271092 542816
rect 146937 542811 147003 542814
rect 271086 542812 271092 542814
rect 271156 542812 271162 542876
rect 322054 542812 322060 542876
rect 322124 542874 322130 542876
rect 358813 542874 358879 542877
rect 322124 542872 358879 542874
rect 322124 542816 358818 542872
rect 358874 542816 358879 542872
rect 322124 542814 358879 542816
rect 322124 542812 322130 542814
rect 358813 542811 358879 542814
rect 363454 542812 363460 542876
rect 363524 542874 363530 542876
rect 391657 542874 391723 542877
rect 363524 542872 391723 542874
rect 363524 542816 391662 542872
rect 391718 542816 391723 542872
rect 363524 542814 391723 542816
rect 363524 542812 363530 542814
rect 391657 542811 391723 542814
rect 197854 542676 197860 542740
rect 197924 542738 197930 542740
rect 336273 542738 336339 542741
rect 197924 542736 336339 542738
rect 197924 542680 336278 542736
rect 336334 542680 336339 542736
rect 197924 542678 336339 542680
rect 197924 542676 197930 542678
rect 336273 542675 336339 542678
rect 367686 542676 367692 542740
rect 367756 542738 367762 542740
rect 380709 542738 380775 542741
rect 367756 542736 380775 542738
rect 367756 542680 380714 542736
rect 380770 542680 380775 542736
rect 367756 542678 380775 542680
rect 367756 542676 367762 542678
rect 380709 542675 380775 542678
rect 113449 542602 113515 542605
rect 137134 542602 137140 542604
rect 113449 542600 137140 542602
rect 113449 542544 113454 542600
rect 113510 542544 137140 542600
rect 113449 542542 137140 542544
rect 113449 542539 113515 542542
rect 137134 542540 137140 542542
rect 137204 542540 137210 542604
rect 149513 542602 149579 542605
rect 166206 542602 166212 542604
rect 149513 542600 166212 542602
rect 149513 542544 149518 542600
rect 149574 542544 166212 542600
rect 149513 542542 166212 542544
rect 149513 542539 149579 542542
rect 166206 542540 166212 542542
rect 166276 542540 166282 542604
rect 210049 542602 210115 542605
rect 222694 542602 222700 542604
rect 210049 542600 222700 542602
rect 210049 542544 210054 542600
rect 210110 542544 222700 542600
rect 210049 542542 222700 542544
rect 210049 542539 210115 542542
rect 222694 542540 222700 542542
rect 222764 542540 222770 542604
rect 242014 542540 242020 542604
rect 242084 542602 242090 542604
rect 251265 542602 251331 542605
rect 242084 542600 251331 542602
rect 242084 542544 251270 542600
rect 251326 542544 251331 542600
rect 242084 542542 251331 542544
rect 242084 542540 242090 542542
rect 251265 542539 251331 542542
rect 266854 542540 266860 542604
rect 266924 542602 266930 542604
rect 353017 542602 353083 542605
rect 266924 542600 353083 542602
rect 266924 542544 353022 542600
rect 353078 542544 353083 542600
rect 266924 542542 353083 542544
rect 266924 542540 266930 542542
rect 353017 542539 353083 542542
rect 353886 542540 353892 542604
rect 353956 542602 353962 542604
rect 366541 542602 366607 542605
rect 353956 542600 366607 542602
rect 353956 542544 366546 542600
rect 366602 542544 366607 542600
rect 353956 542542 366607 542544
rect 353956 542540 353962 542542
rect 366541 542539 366607 542542
rect 389766 542540 389772 542604
rect 389836 542602 389842 542604
rect 396809 542602 396875 542605
rect 389836 542600 396875 542602
rect 389836 542544 396814 542600
rect 396870 542544 396875 542600
rect 389836 542542 396875 542544
rect 389836 542540 389842 542542
rect 396809 542539 396875 542542
rect 138565 542466 138631 542469
rect 152406 542466 152412 542468
rect 138565 542464 152412 542466
rect 138565 542408 138570 542464
rect 138626 542408 152412 542464
rect 138565 542406 152412 542408
rect 138565 542403 138631 542406
rect 152406 542404 152412 542406
rect 152476 542404 152482 542468
rect 161974 542404 161980 542468
rect 162044 542466 162050 542468
rect 177205 542466 177271 542469
rect 162044 542464 177271 542466
rect 162044 542408 177210 542464
rect 177266 542408 177271 542464
rect 162044 542406 177271 542408
rect 162044 542404 162050 542406
rect 177205 542403 177271 542406
rect 190729 542466 190795 542469
rect 208894 542466 208900 542468
rect 190729 542464 208900 542466
rect 190729 542408 190734 542464
rect 190790 542408 208900 542464
rect 190729 542406 208900 542408
rect 190729 542403 190795 542406
rect 208894 542404 208900 542406
rect 208964 542404 208970 542468
rect 231945 542466 232011 542469
rect 237966 542466 237972 542468
rect 231945 542464 237972 542466
rect 231945 542408 231950 542464
rect 232006 542408 237972 542464
rect 231945 542406 237972 542408
rect 231945 542403 232011 542406
rect 237966 542404 237972 542406
rect 238036 542404 238042 542468
rect 250294 542404 250300 542468
rect 250364 542466 250370 542468
rect 257061 542466 257127 542469
rect 250364 542464 257127 542466
rect 250364 542408 257066 542464
rect 257122 542408 257127 542464
rect 250364 542406 257127 542408
rect 250364 542404 250370 542406
rect 257061 542403 257127 542406
rect 215201 541242 215267 541245
rect 215201 541240 238770 541242
rect 215201 541184 215206 541240
rect 215262 541184 238770 541240
rect 215201 541182 238770 541184
rect 215201 541179 215267 541182
rect 238710 541106 238770 541182
rect 304942 541106 304948 541108
rect 238710 541046 304948 541106
rect 304942 541044 304948 541046
rect 305012 541044 305018 541108
rect -960 540684 480 540924
rect 72601 539610 72667 539613
rect 75637 539612 75703 539613
rect 72918 539610 72924 539612
rect 72601 539608 72924 539610
rect 72601 539552 72606 539608
rect 72662 539552 72924 539608
rect 72601 539550 72924 539552
rect 72601 539547 72667 539550
rect 72918 539548 72924 539550
rect 72988 539548 72994 539612
rect 75637 539608 75684 539612
rect 75748 539610 75754 539612
rect 106089 539610 106155 539613
rect 106774 539610 106780 539612
rect 75637 539552 75642 539608
rect 75637 539548 75684 539552
rect 75748 539550 75794 539610
rect 106089 539608 106780 539610
rect 106089 539552 106094 539608
rect 106150 539552 106780 539608
rect 106089 539550 106780 539552
rect 75748 539548 75754 539550
rect 75637 539547 75703 539548
rect 106089 539547 106155 539550
rect 106774 539548 106780 539550
rect 106844 539548 106850 539612
rect 115974 539548 115980 539612
rect 116044 539610 116050 539612
rect 116301 539610 116367 539613
rect 116044 539608 116367 539610
rect 116044 539552 116306 539608
rect 116362 539552 116367 539608
rect 116044 539550 116367 539552
rect 116044 539548 116050 539550
rect 116301 539547 116367 539550
rect 119521 539610 119587 539613
rect 125317 539612 125383 539613
rect 119838 539610 119844 539612
rect 119521 539608 119844 539610
rect 119521 539552 119526 539608
rect 119582 539552 119844 539608
rect 119521 539550 119844 539552
rect 119521 539547 119587 539550
rect 119838 539548 119844 539550
rect 119908 539548 119914 539612
rect 125317 539608 125364 539612
rect 125428 539610 125434 539612
rect 125317 539552 125322 539608
rect 125317 539548 125364 539552
rect 125428 539550 125474 539610
rect 125428 539548 125434 539550
rect 127014 539548 127020 539612
rect 127084 539610 127090 539612
rect 127341 539610 127407 539613
rect 127084 539608 127407 539610
rect 127084 539552 127346 539608
rect 127402 539552 127407 539608
rect 127084 539550 127407 539552
rect 127084 539548 127090 539550
rect 125317 539547 125383 539548
rect 127341 539547 127407 539550
rect 155585 539610 155651 539613
rect 155718 539610 155724 539612
rect 155585 539608 155724 539610
rect 155585 539552 155590 539608
rect 155646 539552 155724 539608
rect 155585 539550 155724 539552
rect 155585 539547 155651 539550
rect 155718 539548 155724 539550
rect 155788 539548 155794 539612
rect 219934 539548 219940 539612
rect 220004 539610 220010 539612
rect 220629 539610 220695 539613
rect 220004 539608 220695 539610
rect 220004 539552 220634 539608
rect 220690 539552 220695 539608
rect 220004 539550 220695 539552
rect 220004 539548 220010 539550
rect 220629 539547 220695 539550
rect 243169 539610 243235 539613
rect 246246 539610 246252 539612
rect 243169 539608 246252 539610
rect 243169 539552 243174 539608
rect 243230 539552 246252 539608
rect 243169 539550 246252 539552
rect 243169 539547 243235 539550
rect 246246 539548 246252 539550
rect 246316 539548 246322 539612
rect 252502 539548 252508 539612
rect 252572 539610 252578 539612
rect 253565 539610 253631 539613
rect 283833 539612 283899 539613
rect 283782 539610 283788 539612
rect 252572 539608 253631 539610
rect 252572 539552 253570 539608
rect 253626 539552 253631 539608
rect 252572 539550 253631 539552
rect 283742 539550 283788 539610
rect 283852 539608 283899 539612
rect 283894 539552 283899 539608
rect 252572 539548 252578 539550
rect 253565 539547 253631 539550
rect 283782 539548 283788 539550
rect 283852 539548 283899 539552
rect 313222 539548 313228 539612
rect 313292 539610 313298 539612
rect 314101 539610 314167 539613
rect 313292 539608 314167 539610
rect 313292 539552 314106 539608
rect 314162 539552 314167 539608
rect 313292 539550 314167 539552
rect 313292 539548 313298 539550
rect 283833 539547 283899 539548
rect 314101 539547 314167 539550
rect 330334 539548 330340 539612
rect 330404 539610 330410 539612
rect 330845 539610 330911 539613
rect 330404 539608 330911 539610
rect 330404 539552 330850 539608
rect 330906 539552 330911 539608
rect 330404 539550 330911 539552
rect 330404 539548 330410 539550
rect 330845 539547 330911 539550
rect 341190 539548 341196 539612
rect 341260 539610 341266 539612
rect 341701 539610 341767 539613
rect 341260 539608 341767 539610
rect 341260 539552 341706 539608
rect 341762 539552 341767 539608
rect 341260 539550 341767 539552
rect 341260 539548 341266 539550
rect 341701 539547 341767 539550
rect 360694 539548 360700 539612
rect 360764 539610 360770 539612
rect 361021 539610 361087 539613
rect 377305 539612 377371 539613
rect 377254 539610 377260 539612
rect 360764 539608 361087 539610
rect 360764 539552 361026 539608
rect 361082 539552 361087 539608
rect 360764 539550 361087 539552
rect 377214 539550 377260 539610
rect 377324 539608 377371 539612
rect 377366 539552 377371 539608
rect 360764 539548 360770 539550
rect 361021 539547 361087 539550
rect 377254 539548 377260 539550
rect 377324 539548 377371 539552
rect 382222 539548 382228 539612
rect 382292 539610 382298 539612
rect 382917 539610 382983 539613
rect 382292 539608 382983 539610
rect 382292 539552 382922 539608
rect 382978 539552 382983 539608
rect 382292 539550 382983 539552
rect 382292 539548 382298 539550
rect 377305 539547 377371 539548
rect 382917 539547 382983 539550
rect 384982 539548 384988 539612
rect 385052 539610 385058 539612
rect 385493 539610 385559 539613
rect 385052 539608 385559 539610
rect 385052 539552 385498 539608
rect 385554 539552 385559 539608
rect 385052 539550 385559 539552
rect 385052 539548 385058 539550
rect 385493 539547 385559 539550
rect 387926 539548 387932 539612
rect 387996 539610 388002 539612
rect 388805 539610 388871 539613
rect 387996 539608 388871 539610
rect 387996 539552 388810 539608
rect 388866 539552 388871 539608
rect 387996 539550 388871 539552
rect 387996 539548 388002 539550
rect 388805 539547 388871 539550
rect 393814 539548 393820 539612
rect 393884 539610 393890 539612
rect 393957 539610 394023 539613
rect 393884 539608 394023 539610
rect 393884 539552 393962 539608
rect 394018 539552 394023 539608
rect 393884 539550 394023 539552
rect 393884 539548 393890 539550
rect 393957 539547 394023 539550
rect 400806 539548 400812 539612
rect 400876 539610 400882 539612
rect 402237 539610 402303 539613
rect 400876 539608 402303 539610
rect 400876 539552 402242 539608
rect 402298 539552 402303 539608
rect 400876 539550 402303 539552
rect 400876 539548 400882 539550
rect 402237 539547 402303 539550
rect 60641 539474 60707 539477
rect 60598 539472 60707 539474
rect 60598 539416 60646 539472
rect 60702 539416 60707 539472
rect 60598 539411 60707 539416
rect 223481 539474 223547 539477
rect 223614 539474 223620 539476
rect 223481 539472 223620 539474
rect 223481 539416 223486 539472
rect 223542 539416 223620 539472
rect 223481 539414 223620 539416
rect 223481 539411 223547 539414
rect 223614 539412 223620 539414
rect 223684 539412 223690 539476
rect 240225 539474 240291 539477
rect 240358 539474 240364 539476
rect 240225 539472 240364 539474
rect 240225 539416 240230 539472
rect 240286 539416 240364 539472
rect 240225 539414 240364 539416
rect 240225 539411 240291 539414
rect 240358 539412 240364 539414
rect 240428 539412 240434 539476
rect 269614 539412 269620 539476
rect 269684 539474 269690 539476
rect 270309 539474 270375 539477
rect 269684 539472 270375 539474
rect 269684 539416 270314 539472
rect 270370 539416 270375 539472
rect 269684 539414 270375 539416
rect 269684 539412 269690 539414
rect 270309 539411 270375 539414
rect 278865 539474 278931 539477
rect 298185 539476 298251 539477
rect 278998 539474 279004 539476
rect 278865 539472 279004 539474
rect 278865 539416 278870 539472
rect 278926 539416 279004 539472
rect 278865 539414 279004 539416
rect 278865 539411 278931 539414
rect 278998 539412 279004 539414
rect 279068 539412 279074 539476
rect 298134 539474 298140 539476
rect 298094 539414 298140 539474
rect 298204 539472 298251 539476
rect 298246 539416 298251 539472
rect 298134 539412 298140 539414
rect 298204 539412 298251 539416
rect 298185 539411 298251 539412
rect 309133 539476 309199 539477
rect 350349 539476 350415 539477
rect 309133 539472 309180 539476
rect 309244 539474 309250 539476
rect 309133 539416 309138 539472
rect 309133 539412 309180 539416
rect 309244 539414 309290 539474
rect 350349 539472 350396 539476
rect 350460 539474 350466 539476
rect 350349 539416 350354 539472
rect 309244 539412 309250 539414
rect 350349 539412 350396 539416
rect 350460 539414 350506 539474
rect 350460 539412 350466 539414
rect 309133 539411 309199 539412
rect 350349 539411 350415 539412
rect 60598 538764 60658 539411
rect 439822 537978 439882 538084
rect 439957 537978 440023 537981
rect 439822 537976 440023 537978
rect 439822 537920 439962 537976
rect 440018 537920 440023 537976
rect 439822 537918 440023 537920
rect 439957 537915 440023 537918
rect 580717 537842 580783 537845
rect 583520 537842 584960 537932
rect 580717 537840 584960 537842
rect 580717 537784 580722 537840
rect 580778 537784 584960 537840
rect 580717 537782 584960 537784
rect 580717 537779 580783 537782
rect 583520 537692 584960 537782
rect 59813 536618 59879 536621
rect 59813 536616 60106 536618
rect 59813 536560 59818 536616
rect 59874 536560 60106 536616
rect 59813 536558 60106 536560
rect 59813 536555 59879 536558
rect 60046 536044 60106 536558
rect 440325 535394 440391 535397
rect 439852 535392 440391 535394
rect 439852 535336 440330 535392
rect 440386 535336 440391 535392
rect 439852 535334 440391 535336
rect 440325 535331 440391 535334
rect 59077 533354 59143 533357
rect 59077 533352 60076 533354
rect 59077 533296 59082 533352
rect 59138 533296 60076 533352
rect 59077 533294 60076 533296
rect 59077 533291 59143 533294
rect 442073 532674 442139 532677
rect 439852 532672 442139 532674
rect 439852 532616 442078 532672
rect 442134 532616 442139 532672
rect 439852 532614 442139 532616
rect 442073 532611 442139 532614
rect 57421 529954 57487 529957
rect 441613 529954 441679 529957
rect 57421 529952 60076 529954
rect 57421 529896 57426 529952
rect 57482 529896 60076 529952
rect 57421 529894 60076 529896
rect 439852 529952 441679 529954
rect 439852 529896 441618 529952
rect 441674 529896 441679 529952
rect 439852 529894 441679 529896
rect 57421 529891 57487 529894
rect 441613 529891 441679 529894
rect -960 527914 480 528004
rect 3233 527914 3299 527917
rect -960 527912 3299 527914
rect -960 527856 3238 527912
rect 3294 527856 3299 527912
rect -960 527854 3299 527856
rect -960 527764 480 527854
rect 3233 527851 3299 527854
rect 57329 527234 57395 527237
rect 57329 527232 60076 527234
rect 57329 527176 57334 527232
rect 57390 527176 60076 527232
rect 57329 527174 60076 527176
rect 57329 527171 57395 527174
rect 440325 526554 440391 526557
rect 439852 526552 440391 526554
rect 439852 526496 440330 526552
rect 440386 526496 440391 526552
rect 439852 526494 440391 526496
rect 440325 526491 440391 526494
rect 57329 524514 57395 524517
rect 580809 524514 580875 524517
rect 583520 524514 584960 524604
rect 57329 524512 60076 524514
rect 57329 524456 57334 524512
rect 57390 524456 60076 524512
rect 57329 524454 60076 524456
rect 580809 524512 584960 524514
rect 580809 524456 580814 524512
rect 580870 524456 584960 524512
rect 580809 524454 584960 524456
rect 57329 524451 57395 524454
rect 580809 524451 580875 524454
rect 583520 524364 584960 524454
rect 442533 523834 442599 523837
rect 439852 523832 442599 523834
rect 439852 523776 442538 523832
rect 442594 523776 442599 523832
rect 439852 523774 442599 523776
rect 442533 523771 442599 523774
rect 57329 521114 57395 521117
rect 440417 521114 440483 521117
rect 57329 521112 60076 521114
rect 57329 521056 57334 521112
rect 57390 521056 60076 521112
rect 57329 521054 60076 521056
rect 439852 521112 440483 521114
rect 439852 521056 440422 521112
rect 440478 521056 440483 521112
rect 439852 521054 440483 521056
rect 57329 521051 57395 521054
rect 440417 521051 440483 521054
rect 57329 518394 57395 518397
rect 57329 518392 60076 518394
rect 57329 518336 57334 518392
rect 57390 518336 60076 518392
rect 57329 518334 60076 518336
rect 57329 518331 57395 518334
rect 442901 517714 442967 517717
rect 439852 517712 442967 517714
rect 439852 517656 442906 517712
rect 442962 517656 442967 517712
rect 439852 517654 442967 517656
rect 442901 517651 442967 517654
rect 57329 515674 57395 515677
rect 57329 515672 60076 515674
rect 57329 515616 57334 515672
rect 57390 515616 60076 515672
rect 57329 515614 60076 515616
rect 57329 515611 57395 515614
rect 442901 514994 442967 514997
rect 439852 514992 442967 514994
rect -960 514858 480 514948
rect 439852 514936 442906 514992
rect 442962 514936 442967 514992
rect 439852 514934 442967 514936
rect 442901 514931 442967 514934
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 57329 512954 57395 512957
rect 57329 512952 60076 512954
rect 57329 512896 57334 512952
rect 57390 512896 60076 512952
rect 57329 512894 60076 512896
rect 57329 512891 57395 512894
rect 442901 512274 442967 512277
rect 439852 512272 442967 512274
rect 439852 512216 442906 512272
rect 442962 512216 442967 512272
rect 439852 512214 442967 512216
rect 442901 512211 442967 512214
rect 580901 511322 580967 511325
rect 583520 511322 584960 511412
rect 580901 511320 584960 511322
rect 580901 511264 580906 511320
rect 580962 511264 584960 511320
rect 580901 511262 584960 511264
rect 580901 511259 580967 511262
rect 583520 511172 584960 511262
rect 57145 509554 57211 509557
rect 442441 509554 442507 509557
rect 57145 509552 60076 509554
rect 57145 509496 57150 509552
rect 57206 509496 60076 509552
rect 57145 509494 60076 509496
rect 439852 509552 442507 509554
rect 439852 509496 442446 509552
rect 442502 509496 442507 509552
rect 439852 509494 442507 509496
rect 57145 509491 57211 509494
rect 442441 509491 442507 509494
rect 56501 506834 56567 506837
rect 56501 506832 60076 506834
rect 56501 506776 56506 506832
rect 56562 506776 60076 506832
rect 56501 506774 60076 506776
rect 56501 506771 56567 506774
rect 442533 506154 442599 506157
rect 439852 506152 442599 506154
rect 439852 506096 442538 506152
rect 442594 506096 442599 506152
rect 439852 506094 442599 506096
rect 442533 506091 442599 506094
rect 57513 504114 57579 504117
rect 57513 504112 60076 504114
rect 57513 504056 57518 504112
rect 57574 504056 60076 504112
rect 57513 504054 60076 504056
rect 57513 504051 57579 504054
rect 442809 503434 442875 503437
rect 439852 503432 442875 503434
rect 439852 503376 442814 503432
rect 442870 503376 442875 503432
rect 439852 503374 442875 503376
rect 442809 503371 442875 503374
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 59169 501394 59235 501397
rect 59169 501392 60076 501394
rect 59169 501336 59174 501392
rect 59230 501336 60076 501392
rect 59169 501334 60076 501336
rect 59169 501331 59235 501334
rect 441797 500714 441863 500717
rect 439852 500712 441863 500714
rect 439852 500656 441802 500712
rect 441858 500656 441863 500712
rect 439852 500654 441863 500656
rect 441797 500651 441863 500654
rect 59353 497994 59419 497997
rect 442533 497994 442599 497997
rect 59353 497992 60076 497994
rect 59353 497936 59358 497992
rect 59414 497936 60076 497992
rect 59353 497934 60076 497936
rect 439852 497992 442599 497994
rect 439852 497936 442538 497992
rect 442594 497936 442599 497992
rect 439852 497934 442599 497936
rect 59353 497931 59419 497934
rect 442533 497931 442599 497934
rect 583520 497844 584960 498084
rect 57605 495274 57671 495277
rect 57605 495272 60076 495274
rect 57605 495216 57610 495272
rect 57666 495216 60076 495272
rect 57605 495214 60076 495216
rect 57605 495211 57671 495214
rect 439865 495138 439931 495141
rect 439822 495136 439931 495138
rect 439822 495080 439870 495136
rect 439926 495080 439931 495136
rect 439822 495075 439931 495080
rect 439822 494564 439882 495075
rect 57605 492554 57671 492557
rect 57605 492552 60076 492554
rect 57605 492496 57610 492552
rect 57666 492496 60076 492552
rect 57605 492494 60076 492496
rect 57605 492491 57671 492494
rect 440417 491874 440483 491877
rect 439852 491872 440483 491874
rect 439852 491816 440422 491872
rect 440478 491816 440483 491872
rect 439852 491814 440483 491816
rect 440417 491811 440483 491814
rect 57605 489154 57671 489157
rect 57605 489152 60076 489154
rect 57605 489096 57610 489152
rect 57666 489096 60076 489152
rect 57605 489094 60076 489096
rect 57605 489091 57671 489094
rect -960 488596 480 488836
rect 439454 488612 439514 489124
rect 439446 488548 439452 488612
rect 439516 488548 439522 488612
rect 442717 486434 442783 486437
rect 439852 486432 442783 486434
rect 60598 485892 60658 486404
rect 439852 486376 442722 486432
rect 442778 486376 442783 486432
rect 439852 486374 442783 486376
rect 442717 486371 442783 486374
rect 60590 485828 60596 485892
rect 60660 485828 60666 485892
rect 580809 484666 580875 484669
rect 583520 484666 584960 484756
rect 580809 484664 584960 484666
rect 580809 484608 580814 484664
rect 580870 484608 584960 484664
rect 580809 484606 584960 484608
rect 580809 484603 580875 484606
rect 583520 484516 584960 484606
rect 57789 483714 57855 483717
rect 57789 483712 60076 483714
rect 57789 483656 57794 483712
rect 57850 483656 60076 483712
rect 57789 483654 60076 483656
rect 57789 483651 57855 483654
rect 441797 483034 441863 483037
rect 439852 483032 441863 483034
rect 439852 482976 441802 483032
rect 441858 482976 441863 483032
rect 439852 482974 441863 482976
rect 441797 482971 441863 482974
rect 57605 480994 57671 480997
rect 57605 480992 60076 480994
rect 57605 480936 57610 480992
rect 57666 480936 60076 480992
rect 57605 480934 60076 480936
rect 57605 480931 57671 480934
rect 442901 480314 442967 480317
rect 439852 480312 442967 480314
rect 439852 480256 442906 480312
rect 442962 480256 442967 480312
rect 439852 480254 442967 480256
rect 442901 480251 442967 480254
rect 57053 477594 57119 477597
rect 441889 477594 441955 477597
rect 57053 477592 60076 477594
rect 57053 477536 57058 477592
rect 57114 477536 60076 477592
rect 57053 477534 60076 477536
rect 439852 477592 441955 477594
rect 439852 477536 441894 477592
rect 441950 477536 441955 477592
rect 439852 477534 441955 477536
rect 57053 477531 57119 477534
rect 441889 477531 441955 477534
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 57605 474874 57671 474877
rect 57605 474872 60076 474874
rect 57605 474816 57610 474872
rect 57666 474816 60076 474872
rect 57605 474814 60076 474816
rect 57605 474811 57671 474814
rect 442901 474194 442967 474197
rect 439852 474192 442967 474194
rect 439852 474136 442906 474192
rect 442962 474136 442967 474192
rect 439852 474134 442967 474136
rect 442901 474131 442967 474134
rect 58985 472154 59051 472157
rect 58985 472152 60076 472154
rect 58985 472096 58990 472152
rect 59046 472096 60076 472152
rect 58985 472094 60076 472096
rect 58985 472091 59051 472094
rect 442901 471474 442967 471477
rect 439852 471472 442967 471474
rect 439852 471416 442906 471472
rect 442962 471416 442967 471472
rect 439852 471414 442967 471416
rect 442901 471411 442967 471414
rect 580441 471474 580507 471477
rect 583520 471474 584960 471564
rect 580441 471472 584960 471474
rect 580441 471416 580446 471472
rect 580502 471416 584960 471472
rect 580441 471414 584960 471416
rect 580441 471411 580507 471414
rect 583520 471324 584960 471414
rect 57605 469434 57671 469437
rect 57605 469432 60076 469434
rect 57605 469376 57610 469432
rect 57666 469376 60076 469432
rect 57605 469374 60076 469376
rect 57605 469371 57671 469374
rect 442901 468754 442967 468757
rect 439852 468752 442967 468754
rect 439852 468696 442906 468752
rect 442962 468696 442967 468752
rect 439852 468694 442967 468696
rect 442901 468691 442967 468694
rect 56869 466034 56935 466037
rect 442809 466034 442875 466037
rect 56869 466032 60076 466034
rect 56869 465976 56874 466032
rect 56930 465976 60076 466032
rect 56869 465974 60076 465976
rect 439852 466032 442875 466034
rect 439852 465976 442814 466032
rect 442870 465976 442875 466032
rect 439852 465974 442875 465976
rect 56869 465971 56935 465974
rect 442809 465971 442875 465974
rect 57605 463314 57671 463317
rect 57605 463312 60076 463314
rect 57605 463256 57610 463312
rect 57666 463256 60076 463312
rect 57605 463254 60076 463256
rect 57605 463251 57671 463254
rect -960 462634 480 462724
rect 442901 462634 442967 462637
rect -960 462574 6930 462634
rect 439852 462632 442967 462634
rect 439852 462576 442906 462632
rect 442962 462576 442967 462632
rect 439852 462574 442967 462576
rect -960 462484 480 462574
rect 6870 462362 6930 462574
rect 442901 462571 442967 462574
rect 33726 462362 33732 462364
rect 6870 462302 33732 462362
rect 33726 462300 33732 462302
rect 33796 462300 33802 462364
rect 57605 460594 57671 460597
rect 57605 460592 60076 460594
rect 57605 460536 57610 460592
rect 57666 460536 60076 460592
rect 57605 460534 60076 460536
rect 57605 460531 57671 460534
rect 442901 459914 442967 459917
rect 439852 459912 442967 459914
rect 439852 459856 442906 459912
rect 442962 459856 442967 459912
rect 439852 459854 442967 459856
rect 442901 459851 442967 459854
rect 580441 458146 580507 458149
rect 583520 458146 584960 458236
rect 580441 458144 584960 458146
rect 580441 458088 580446 458144
rect 580502 458088 584960 458144
rect 580441 458086 584960 458088
rect 580441 458083 580507 458086
rect 583520 457996 584960 458086
rect 57605 457874 57671 457877
rect 57605 457872 60076 457874
rect 57605 457816 57610 457872
rect 57666 457816 60076 457872
rect 57605 457814 60076 457816
rect 57605 457811 57671 457814
rect 442901 457194 442967 457197
rect 439852 457192 442967 457194
rect 439852 457136 442906 457192
rect 442962 457136 442967 457192
rect 439852 457134 442967 457136
rect 442901 457131 442967 457134
rect 57605 454474 57671 454477
rect 442901 454474 442967 454477
rect 57605 454472 60076 454474
rect 57605 454416 57610 454472
rect 57666 454416 60076 454472
rect 57605 454414 60076 454416
rect 439852 454472 442967 454474
rect 439852 454416 442906 454472
rect 442962 454416 442967 454472
rect 439852 454414 442967 454416
rect 57605 454411 57671 454414
rect 442901 454411 442967 454414
rect 57605 451754 57671 451757
rect 57605 451752 60076 451754
rect 57605 451696 57610 451752
rect 57666 451696 60076 451752
rect 57605 451694 60076 451696
rect 57605 451691 57671 451694
rect 440693 451074 440759 451077
rect 439852 451072 440759 451074
rect 439852 451016 440698 451072
rect 440754 451016 440759 451072
rect 439852 451014 440759 451016
rect 440693 451011 440759 451014
rect -960 449578 480 449668
rect 3969 449578 4035 449581
rect -960 449576 4035 449578
rect -960 449520 3974 449576
rect 4030 449520 4035 449576
rect -960 449518 4035 449520
rect -960 449428 480 449518
rect 3969 449515 4035 449518
rect 57789 449034 57855 449037
rect 57789 449032 60076 449034
rect 57789 448976 57794 449032
rect 57850 448976 60076 449032
rect 57789 448974 60076 448976
rect 57789 448971 57855 448974
rect 442901 448354 442967 448357
rect 439852 448352 442967 448354
rect 439852 448296 442906 448352
rect 442962 448296 442967 448352
rect 439852 448294 442967 448296
rect 442901 448291 442967 448294
rect 439497 445906 439563 445909
rect 439454 445904 439563 445906
rect 439454 445848 439502 445904
rect 439558 445848 439563 445904
rect 439454 445843 439563 445848
rect 57053 445634 57119 445637
rect 57053 445632 60076 445634
rect 57053 445576 57058 445632
rect 57114 445576 60076 445632
rect 439454 445604 439514 445843
rect 57053 445574 60076 445576
rect 57053 445571 57119 445574
rect 583520 444668 584960 444908
rect 56409 442914 56475 442917
rect 56409 442912 60076 442914
rect 56409 442856 56414 442912
rect 56470 442856 60076 442912
rect 56409 442854 60076 442856
rect 56409 442851 56475 442854
rect 442349 442234 442415 442237
rect 439852 442232 442415 442234
rect 439852 442176 442354 442232
rect 442410 442176 442415 442232
rect 439852 442174 442415 442176
rect 442349 442171 442415 442174
rect 56317 440194 56383 440197
rect 56317 440192 60076 440194
rect 56317 440136 56322 440192
rect 56378 440136 60076 440192
rect 56317 440134 60076 440136
rect 56317 440131 56383 440134
rect 439454 438973 439514 439484
rect 439454 438968 439563 438973
rect 439454 438912 439502 438968
rect 439558 438912 439563 438968
rect 439454 438910 439563 438912
rect 439497 438907 439563 438910
rect 57605 437474 57671 437477
rect 57605 437472 60076 437474
rect 57605 437416 57610 437472
rect 57666 437416 60076 437472
rect 57605 437414 60076 437416
rect 57605 437411 57671 437414
rect 442717 436794 442783 436797
rect 439852 436792 442783 436794
rect -960 436508 480 436748
rect 439852 436736 442722 436792
rect 442778 436736 442783 436792
rect 439852 436734 442783 436736
rect 442717 436731 442783 436734
rect 57605 434074 57671 434077
rect 57605 434072 60076 434074
rect 57605 434016 57610 434072
rect 57666 434016 60076 434072
rect 57605 434014 60076 434016
rect 57605 434011 57671 434014
rect 439454 433532 439514 434044
rect 439446 433468 439452 433532
rect 439516 433468 439522 433532
rect 579981 431626 580047 431629
rect 583520 431626 584960 431716
rect 579981 431624 584960 431626
rect 579981 431568 579986 431624
rect 580042 431568 584960 431624
rect 579981 431566 584960 431568
rect 579981 431563 580047 431566
rect 583520 431476 584960 431566
rect 57605 431354 57671 431357
rect 57605 431352 60076 431354
rect 57605 431296 57610 431352
rect 57666 431296 60076 431352
rect 57605 431294 60076 431296
rect 57605 431291 57671 431294
rect 442901 430674 442967 430677
rect 439852 430672 442967 430674
rect 439852 430616 442906 430672
rect 442962 430616 442967 430672
rect 439852 430614 442967 430616
rect 442901 430611 442967 430614
rect 57605 428634 57671 428637
rect 57605 428632 60076 428634
rect 57605 428576 57610 428632
rect 57666 428576 60076 428632
rect 57605 428574 60076 428576
rect 57605 428571 57671 428574
rect 440785 427954 440851 427957
rect 439852 427952 440851 427954
rect 439852 427896 440790 427952
rect 440846 427896 440851 427952
rect 439852 427894 440851 427896
rect 440785 427891 440851 427894
rect 59445 425914 59511 425917
rect 59445 425912 60076 425914
rect 59445 425856 59450 425912
rect 59506 425856 60076 425912
rect 59445 425854 60076 425856
rect 59445 425851 59511 425854
rect 439262 425716 439268 425780
rect 439332 425716 439338 425780
rect 439270 425204 439330 425716
rect -960 423602 480 423692
rect 3693 423602 3759 423605
rect -960 423600 3759 423602
rect -960 423544 3698 423600
rect 3754 423544 3759 423600
rect -960 423542 3759 423544
rect -960 423452 480 423542
rect 3693 423539 3759 423542
rect 57605 422514 57671 422517
rect 442901 422514 442967 422517
rect 57605 422512 60076 422514
rect 57605 422456 57610 422512
rect 57666 422456 60076 422512
rect 57605 422454 60076 422456
rect 439852 422512 442967 422514
rect 439852 422456 442906 422512
rect 442962 422456 442967 422512
rect 439852 422454 442967 422456
rect 57605 422451 57671 422454
rect 442901 422451 442967 422454
rect 57605 419794 57671 419797
rect 57605 419792 60076 419794
rect 57605 419736 57610 419792
rect 57666 419736 60076 419792
rect 57605 419734 60076 419736
rect 57605 419731 57671 419734
rect 442533 419114 442599 419117
rect 439852 419112 442599 419114
rect 439852 419056 442538 419112
rect 442594 419056 442599 419112
rect 439852 419054 442599 419056
rect 442533 419051 442599 419054
rect 453246 418236 453252 418300
rect 453316 418298 453322 418300
rect 583520 418298 584960 418388
rect 453316 418238 584960 418298
rect 453316 418236 453322 418238
rect 583520 418148 584960 418238
rect 57605 417074 57671 417077
rect 57605 417072 60076 417074
rect 57605 417016 57610 417072
rect 57666 417016 60076 417072
rect 57605 417014 60076 417016
rect 57605 417011 57671 417014
rect 442717 416394 442783 416397
rect 439852 416392 442783 416394
rect 439852 416336 442722 416392
rect 442778 416336 442783 416392
rect 439852 416334 442783 416336
rect 442717 416331 442783 416334
rect 57605 413674 57671 413677
rect 443177 413674 443243 413677
rect 57605 413672 60076 413674
rect 57605 413616 57610 413672
rect 57666 413616 60076 413672
rect 57605 413614 60076 413616
rect 439852 413672 443243 413674
rect 439852 413616 443182 413672
rect 443238 413616 443243 413672
rect 439852 413614 443243 413616
rect 57605 413611 57671 413614
rect 443177 413611 443243 413614
rect 57513 410954 57579 410957
rect 57513 410952 60076 410954
rect 57513 410896 57518 410952
rect 57574 410896 60076 410952
rect 57513 410894 60076 410896
rect 57513 410891 57579 410894
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 442533 410274 442599 410277
rect 439852 410272 442599 410274
rect 439852 410216 442538 410272
rect 442594 410216 442599 410272
rect 439852 410214 442599 410216
rect 442533 410211 442599 410214
rect 56225 408234 56291 408237
rect 56225 408232 60076 408234
rect 56225 408176 56230 408232
rect 56286 408176 60076 408232
rect 56225 408174 60076 408176
rect 56225 408171 56291 408174
rect 441981 407554 442047 407557
rect 439852 407552 442047 407554
rect 439852 407496 441986 407552
rect 442042 407496 442047 407552
rect 439852 407494 442047 407496
rect 441981 407491 442047 407494
rect 58893 405514 58959 405517
rect 58893 405512 60076 405514
rect 58893 405456 58898 405512
rect 58954 405456 60076 405512
rect 58893 405454 60076 405456
rect 58893 405451 58959 405454
rect 583520 404970 584960 405060
rect 583342 404910 584960 404970
rect 442533 404834 442599 404837
rect 439852 404832 442599 404834
rect 439852 404776 442538 404832
rect 442594 404776 442599 404832
rect 439852 404774 442599 404776
rect 583342 404834 583402 404910
rect 583520 404834 584960 404910
rect 583342 404820 584960 404834
rect 583342 404774 583586 404820
rect 442533 404771 442599 404774
rect 450486 404364 450492 404428
rect 450556 404426 450562 404428
rect 583526 404426 583586 404774
rect 450556 404366 583586 404426
rect 450556 404364 450562 404366
rect 57513 402114 57579 402117
rect 442073 402114 442139 402117
rect 57513 402112 60076 402114
rect 57513 402056 57518 402112
rect 57574 402056 60076 402112
rect 57513 402054 60076 402056
rect 439852 402112 442139 402114
rect 439852 402056 442078 402112
rect 442134 402056 442139 402112
rect 439852 402054 442139 402056
rect 57513 402051 57579 402054
rect 442073 402051 442139 402054
rect 57513 399394 57579 399397
rect 57513 399392 60076 399394
rect 57513 399336 57518 399392
rect 57574 399336 60076 399392
rect 57513 399334 60076 399336
rect 57513 399331 57579 399334
rect 3601 398714 3667 398717
rect 21214 398714 21220 398716
rect 3601 398712 21220 398714
rect 3601 398656 3606 398712
rect 3662 398656 21220 398712
rect 3601 398654 21220 398656
rect 3601 398651 3667 398654
rect 21214 398652 21220 398654
rect 21284 398652 21290 398716
rect 439454 398172 439514 398684
rect 439446 398108 439452 398172
rect 439516 398108 439522 398172
rect -960 397490 480 397580
rect 3601 397490 3667 397493
rect -960 397488 3667 397490
rect -960 397432 3606 397488
rect 3662 397432 3667 397488
rect -960 397430 3667 397432
rect -960 397340 480 397430
rect 3601 397427 3667 397430
rect 57513 396674 57579 396677
rect 57513 396672 60076 396674
rect 57513 396616 57518 396672
rect 57574 396616 60076 396672
rect 57513 396614 60076 396616
rect 57513 396611 57579 396614
rect 442901 395994 442967 395997
rect 439852 395992 442967 395994
rect 439852 395936 442906 395992
rect 442962 395936 442967 395992
rect 439852 395934 442967 395936
rect 442901 395931 442967 395934
rect 57513 393954 57579 393957
rect 57513 393952 60076 393954
rect 57513 393896 57518 393952
rect 57574 393896 60076 393952
rect 57513 393894 60076 393896
rect 57513 393891 57579 393894
rect 439454 392732 439514 393244
rect 439446 392668 439452 392732
rect 439516 392668 439522 392732
rect 583520 391628 584960 391868
rect 57513 390554 57579 390557
rect 442257 390554 442323 390557
rect 57513 390552 60076 390554
rect 57513 390496 57518 390552
rect 57574 390496 60076 390552
rect 57513 390494 60076 390496
rect 439852 390552 442323 390554
rect 439852 390496 442262 390552
rect 442318 390496 442323 390552
rect 439852 390494 442323 390496
rect 57513 390491 57579 390494
rect 442257 390491 442323 390494
rect 57513 387834 57579 387837
rect 57513 387832 60076 387834
rect 57513 387776 57518 387832
rect 57574 387776 60076 387832
rect 57513 387774 60076 387776
rect 57513 387771 57579 387774
rect 439773 387698 439839 387701
rect 439773 387696 439882 387698
rect 439773 387640 439778 387696
rect 439834 387640 439882 387696
rect 439773 387635 439882 387640
rect 439822 387124 439882 387635
rect 57513 385114 57579 385117
rect 57513 385112 60076 385114
rect 57513 385056 57518 385112
rect 57574 385056 60076 385112
rect 57513 385054 60076 385056
rect 57513 385051 57579 385054
rect -960 384284 480 384524
rect 440785 384434 440851 384437
rect 439852 384432 440851 384434
rect 439852 384376 440790 384432
rect 440846 384376 440851 384432
rect 439852 384374 440851 384376
rect 440785 384371 440851 384374
rect 57513 381714 57579 381717
rect 442901 381714 442967 381717
rect 57513 381712 60076 381714
rect 57513 381656 57518 381712
rect 57574 381656 60076 381712
rect 57513 381654 60076 381656
rect 439852 381712 442967 381714
rect 439852 381656 442906 381712
rect 442962 381656 442967 381712
rect 439852 381654 442967 381656
rect 57513 381651 57579 381654
rect 442901 381651 442967 381654
rect 57513 378994 57579 378997
rect 442901 378994 442967 378997
rect 57513 378992 60076 378994
rect 57513 378936 57518 378992
rect 57574 378936 60076 378992
rect 57513 378934 60076 378936
rect 439852 378992 442967 378994
rect 439852 378936 442906 378992
rect 442962 378936 442967 378992
rect 439852 378934 442967 378936
rect 57513 378931 57579 378934
rect 442901 378931 442967 378934
rect 583520 378450 584960 378540
rect 567150 378390 584960 378450
rect 500166 378116 500172 378180
rect 500236 378178 500242 378180
rect 567150 378178 567210 378390
rect 583520 378300 584960 378390
rect 500236 378118 567210 378178
rect 500236 378116 500242 378118
rect 58801 376274 58867 376277
rect 58801 376272 60076 376274
rect 58801 376216 58806 376272
rect 58862 376216 60076 376272
rect 58801 376214 60076 376216
rect 58801 376211 58867 376214
rect 442901 375594 442967 375597
rect 439852 375592 442967 375594
rect 439852 375536 442906 375592
rect 442962 375536 442967 375592
rect 439852 375534 442967 375536
rect 442901 375531 442967 375534
rect 57513 373554 57579 373557
rect 57513 373552 60076 373554
rect 57513 373496 57518 373552
rect 57574 373496 60076 373552
rect 57513 373494 60076 373496
rect 57513 373491 57579 373494
rect 442901 372874 442967 372877
rect 439852 372872 442967 372874
rect 439852 372816 442906 372872
rect 442962 372816 442967 372872
rect 439852 372814 442967 372816
rect 442901 372811 442967 372814
rect -960 371378 480 371468
rect 3601 371378 3667 371381
rect -960 371376 3667 371378
rect -960 371320 3606 371376
rect 3662 371320 3667 371376
rect -960 371318 3667 371320
rect -960 371228 480 371318
rect 3601 371315 3667 371318
rect 60590 370636 60596 370700
rect 60660 370636 60666 370700
rect 60598 370124 60658 370636
rect 442165 370154 442231 370157
rect 439852 370152 442231 370154
rect 439852 370096 442170 370152
rect 442226 370096 442231 370152
rect 439852 370094 442231 370096
rect 442165 370091 442231 370094
rect 56869 367434 56935 367437
rect 56869 367432 60076 367434
rect 56869 367376 56874 367432
rect 56930 367376 60076 367432
rect 56869 367374 60076 367376
rect 56869 367371 56935 367374
rect 442901 366754 442967 366757
rect 439852 366752 442967 366754
rect 439852 366696 442906 366752
rect 442962 366696 442967 366752
rect 439852 366694 442967 366696
rect 442901 366691 442967 366694
rect 579981 365122 580047 365125
rect 583520 365122 584960 365212
rect 579981 365120 584960 365122
rect 579981 365064 579986 365120
rect 580042 365064 584960 365120
rect 579981 365062 584960 365064
rect 579981 365059 580047 365062
rect 583520 364972 584960 365062
rect 56869 364714 56935 364717
rect 56869 364712 60076 364714
rect 56869 364656 56874 364712
rect 56930 364656 60076 364712
rect 56869 364654 60076 364656
rect 56869 364651 56935 364654
rect 443085 364034 443151 364037
rect 439852 364032 443151 364034
rect 439852 363976 443090 364032
rect 443146 363976 443151 364032
rect 439852 363974 443151 363976
rect 443085 363971 443151 363974
rect 57513 361994 57579 361997
rect 57513 361992 60076 361994
rect 57513 361936 57518 361992
rect 57574 361936 60076 361992
rect 57513 361934 60076 361936
rect 57513 361931 57579 361934
rect 442625 361314 442691 361317
rect 439852 361312 442691 361314
rect 439852 361256 442630 361312
rect 442686 361256 442691 361312
rect 439852 361254 442691 361256
rect 442625 361251 442691 361254
rect 57513 358594 57579 358597
rect 442717 358594 442783 358597
rect 57513 358592 60076 358594
rect -960 358458 480 358548
rect 57513 358536 57518 358592
rect 57574 358536 60076 358592
rect 57513 358534 60076 358536
rect 439852 358592 442783 358594
rect 439852 358536 442722 358592
rect 442778 358536 442783 358592
rect 439852 358534 442783 358536
rect 57513 358531 57579 358534
rect 442717 358531 442783 358534
rect 3693 358458 3759 358461
rect -960 358456 3759 358458
rect -960 358400 3698 358456
rect 3754 358400 3759 358456
rect -960 358398 3759 358400
rect -960 358308 480 358398
rect 3693 358395 3759 358398
rect 56041 355874 56107 355877
rect 56041 355872 60076 355874
rect 56041 355816 56046 355872
rect 56102 355816 60076 355872
rect 56041 355814 60076 355816
rect 56041 355811 56107 355814
rect 442901 355194 442967 355197
rect 439852 355192 442967 355194
rect 439852 355136 442906 355192
rect 442962 355136 442967 355192
rect 439852 355134 442967 355136
rect 442901 355131 442967 355134
rect 57513 353154 57579 353157
rect 57513 353152 60076 353154
rect 57513 353096 57518 353152
rect 57574 353096 60076 353152
rect 57513 353094 60076 353096
rect 57513 353091 57579 353094
rect 442901 352474 442967 352477
rect 439852 352472 442967 352474
rect 439852 352416 442906 352472
rect 442962 352416 442967 352472
rect 439852 352414 442967 352416
rect 442901 352411 442967 352414
rect 580073 351930 580139 351933
rect 583520 351930 584960 352020
rect 580073 351928 584960 351930
rect 580073 351872 580078 351928
rect 580134 351872 584960 351928
rect 580073 351870 584960 351872
rect 580073 351867 580139 351870
rect 583520 351780 584960 351870
rect 56869 350434 56935 350437
rect 56869 350432 60076 350434
rect 56869 350376 56874 350432
rect 56930 350376 60076 350432
rect 56869 350374 60076 350376
rect 56869 350371 56935 350374
rect 442717 349754 442783 349757
rect 439852 349752 442783 349754
rect 439852 349696 442722 349752
rect 442778 349696 442783 349752
rect 439852 349694 442783 349696
rect 442717 349691 442783 349694
rect 439446 347244 439452 347308
rect 439516 347244 439522 347308
rect 57513 347034 57579 347037
rect 57513 347032 60076 347034
rect 57513 346976 57518 347032
rect 57574 346976 60076 347032
rect 439454 347004 439514 347244
rect 57513 346974 60076 346976
rect 57513 346971 57579 346974
rect -960 345402 480 345492
rect 3785 345402 3851 345405
rect -960 345400 3851 345402
rect -960 345344 3790 345400
rect 3846 345344 3851 345400
rect -960 345342 3851 345344
rect -960 345252 480 345342
rect 3785 345339 3851 345342
rect 60598 343772 60658 344284
rect 60590 343708 60596 343772
rect 60660 343708 60666 343772
rect 442901 343634 442967 343637
rect 439852 343632 442967 343634
rect 439852 343576 442906 343632
rect 442962 343576 442967 343632
rect 439852 343574 442967 343576
rect 442901 343571 442967 343574
rect 57513 341594 57579 341597
rect 57513 341592 60076 341594
rect 57513 341536 57518 341592
rect 57574 341536 60076 341592
rect 57513 341534 60076 341536
rect 57513 341531 57579 341534
rect 442901 340914 442967 340917
rect 439852 340912 442967 340914
rect 439852 340856 442906 340912
rect 442962 340856 442967 340912
rect 439852 340854 442967 340856
rect 442901 340851 442967 340854
rect 583520 338452 584960 338692
rect 57513 338194 57579 338197
rect 442901 338194 442967 338197
rect 57513 338192 60076 338194
rect 57513 338136 57518 338192
rect 57574 338136 60076 338192
rect 57513 338134 60076 338136
rect 439852 338192 442967 338194
rect 439852 338136 442906 338192
rect 442962 338136 442967 338192
rect 439852 338134 442967 338136
rect 57513 338131 57579 338134
rect 442901 338131 442967 338134
rect 55949 335474 56015 335477
rect 55949 335472 60076 335474
rect 55949 335416 55954 335472
rect 56010 335416 60076 335472
rect 55949 335414 60076 335416
rect 55949 335411 56015 335414
rect 442717 334794 442783 334797
rect 439852 334792 442783 334794
rect 439852 334736 442722 334792
rect 442778 334736 442783 334792
rect 439852 334734 442783 334736
rect 442717 334731 442783 334734
rect 57881 332754 57947 332757
rect 57881 332752 60076 332754
rect 57881 332696 57886 332752
rect 57942 332696 60076 332752
rect 57881 332694 60076 332696
rect 57881 332691 57947 332694
rect -960 332196 480 332436
rect 442901 332074 442967 332077
rect 439852 332072 442967 332074
rect 439852 332016 442906 332072
rect 442962 332016 442967 332072
rect 439852 332014 442967 332016
rect 442901 332011 442967 332014
rect 57513 330034 57579 330037
rect 57513 330032 60076 330034
rect 57513 329976 57518 330032
rect 57574 329976 60076 330032
rect 57513 329974 60076 329976
rect 57513 329971 57579 329974
rect 442901 329354 442967 329357
rect 439852 329352 442967 329354
rect 439852 329296 442906 329352
rect 442962 329296 442967 329352
rect 439852 329294 442967 329296
rect 442901 329291 442967 329294
rect 56133 326634 56199 326637
rect 442533 326634 442599 326637
rect 56133 326632 60076 326634
rect 56133 326576 56138 326632
rect 56194 326576 60076 326632
rect 56133 326574 60076 326576
rect 439852 326632 442599 326634
rect 439852 326576 442538 326632
rect 442594 326576 442599 326632
rect 439852 326574 442599 326576
rect 56133 326571 56199 326574
rect 442533 326571 442599 326574
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 57329 323914 57395 323917
rect 57329 323912 60076 323914
rect 57329 323856 57334 323912
rect 57390 323856 60076 323912
rect 57329 323854 60076 323856
rect 57329 323851 57395 323854
rect 442533 323234 442599 323237
rect 439852 323232 442599 323234
rect 439852 323176 442538 323232
rect 442594 323176 442599 323232
rect 439852 323174 442599 323176
rect 442533 323171 442599 323174
rect 57973 321194 58039 321197
rect 57973 321192 60076 321194
rect 57973 321136 57978 321192
rect 58034 321136 60076 321192
rect 57973 321134 60076 321136
rect 57973 321131 58039 321134
rect 442901 320514 442967 320517
rect 439852 320512 442967 320514
rect 439852 320456 442906 320512
rect 442962 320456 442967 320512
rect 439852 320454 442967 320456
rect 442901 320451 442967 320454
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 59537 318474 59603 318477
rect 59537 318472 60076 318474
rect 59537 318416 59542 318472
rect 59598 318416 60076 318472
rect 59537 318414 60076 318416
rect 59537 318411 59603 318414
rect 442901 317794 442967 317797
rect 439852 317792 442967 317794
rect 439852 317736 442906 317792
rect 442962 317736 442967 317792
rect 439852 317734 442967 317736
rect 442901 317731 442967 317734
rect 56869 315074 56935 315077
rect 442257 315074 442323 315077
rect 56869 315072 60076 315074
rect 56869 315016 56874 315072
rect 56930 315016 60076 315072
rect 56869 315014 60076 315016
rect 439852 315072 442323 315074
rect 439852 315016 442262 315072
rect 442318 315016 442323 315072
rect 439852 315014 442323 315016
rect 56869 315011 56935 315014
rect 442257 315011 442323 315014
rect 57329 312354 57395 312357
rect 57329 312352 60076 312354
rect 57329 312296 57334 312352
rect 57390 312296 60076 312352
rect 57329 312294 60076 312296
rect 57329 312291 57395 312294
rect 583520 312082 584960 312172
rect 567150 312022 584960 312082
rect 471094 311884 471100 311948
rect 471164 311946 471170 311948
rect 567150 311946 567210 312022
rect 471164 311886 567210 311946
rect 583520 311932 584960 312022
rect 471164 311884 471170 311886
rect 442717 311674 442783 311677
rect 439852 311672 442783 311674
rect 439852 311616 442722 311672
rect 442778 311616 442783 311672
rect 439852 311614 442783 311616
rect 442717 311611 442783 311614
rect 57329 309634 57395 309637
rect 57329 309632 60076 309634
rect 57329 309576 57334 309632
rect 57390 309576 60076 309632
rect 57329 309574 60076 309576
rect 57329 309571 57395 309574
rect 442901 308954 442967 308957
rect 439852 308952 442967 308954
rect 439852 308896 442906 308952
rect 442962 308896 442967 308952
rect 439852 308894 442967 308896
rect 442901 308891 442967 308894
rect 35014 306370 35020 306372
rect -960 306234 480 306324
rect 6870 306310 35020 306370
rect 6870 306234 6930 306310
rect 35014 306308 35020 306310
rect 35084 306308 35090 306372
rect -960 306174 6930 306234
rect 59629 306234 59695 306237
rect 440877 306234 440943 306237
rect 59629 306232 60076 306234
rect 59629 306176 59634 306232
rect 59690 306176 60076 306232
rect 59629 306174 60076 306176
rect 439852 306232 440943 306234
rect 439852 306176 440882 306232
rect 440938 306176 440943 306232
rect 439852 306174 440943 306176
rect -960 306084 480 306174
rect 59629 306171 59695 306174
rect 440877 306171 440943 306174
rect 60598 303380 60658 303484
rect 60590 303316 60596 303380
rect 60660 303316 60666 303380
rect 442441 302834 442507 302837
rect 439852 302832 442507 302834
rect 439852 302776 442446 302832
rect 442502 302776 442507 302832
rect 439852 302774 442507 302776
rect 442441 302771 442507 302774
rect 439446 302092 439452 302156
rect 439516 302154 439522 302156
rect 449934 302154 449940 302156
rect 439516 302094 449940 302154
rect 439516 302092 439522 302094
rect 449934 302092 449940 302094
rect 450004 302092 450010 302156
rect 57329 300794 57395 300797
rect 57329 300792 60076 300794
rect 57329 300736 57334 300792
rect 57390 300736 60076 300792
rect 57329 300734 60076 300736
rect 57329 300731 57395 300734
rect 440969 300114 441035 300117
rect 439852 300112 441035 300114
rect 439852 300056 440974 300112
rect 441030 300056 441035 300112
rect 439852 300054 441035 300056
rect 440969 300051 441035 300054
rect 583520 298754 584960 298844
rect 583342 298694 584960 298754
rect 583342 298618 583402 298694
rect 583520 298618 584960 298694
rect 583342 298604 584960 298618
rect 583342 298558 583586 298604
rect 449934 298148 449940 298212
rect 450004 298210 450010 298212
rect 583526 298210 583586 298558
rect 450004 298150 583586 298210
rect 450004 298148 450010 298150
rect 57329 298074 57395 298077
rect 57329 298072 60076 298074
rect 57329 298016 57334 298072
rect 57390 298016 60076 298072
rect 57329 298014 60076 298016
rect 57329 298011 57395 298014
rect 442901 297394 442967 297397
rect 439852 297392 442967 297394
rect 439852 297336 442906 297392
rect 442962 297336 442967 297392
rect 439852 297334 442967 297336
rect 442901 297331 442967 297334
rect 57881 294674 57947 294677
rect 442441 294674 442507 294677
rect 57881 294672 60076 294674
rect 57881 294616 57886 294672
rect 57942 294616 60076 294672
rect 57881 294614 60076 294616
rect 439852 294672 442507 294674
rect 439852 294616 442446 294672
rect 442502 294616 442507 294672
rect 439852 294614 442507 294616
rect 57881 294611 57947 294614
rect 442441 294611 442507 294614
rect -960 293178 480 293268
rect 3969 293178 4035 293181
rect -960 293176 4035 293178
rect -960 293120 3974 293176
rect 4030 293120 4035 293176
rect -960 293118 4035 293120
rect -960 293028 480 293118
rect 3969 293115 4035 293118
rect 57053 291954 57119 291957
rect 57053 291952 60076 291954
rect 57053 291896 57058 291952
rect 57114 291896 60076 291952
rect 57053 291894 60076 291896
rect 57053 291891 57119 291894
rect 442901 291274 442967 291277
rect 439852 291272 442967 291274
rect 439852 291216 442906 291272
rect 442962 291216 442967 291272
rect 439852 291214 442967 291216
rect 442901 291211 442967 291214
rect 57329 289234 57395 289237
rect 57329 289232 60076 289234
rect 57329 289176 57334 289232
rect 57390 289176 60076 289232
rect 57329 289174 60076 289176
rect 57329 289171 57395 289174
rect 442901 288554 442967 288557
rect 439852 288552 442967 288554
rect 439852 288496 442906 288552
rect 442962 288496 442967 288552
rect 439852 288494 442967 288496
rect 442901 288491 442967 288494
rect 58709 286514 58775 286517
rect 58709 286512 60076 286514
rect 58709 286456 58714 286512
rect 58770 286456 60076 286512
rect 58709 286454 60076 286456
rect 58709 286451 58775 286454
rect 442901 285834 442967 285837
rect 439852 285832 442967 285834
rect 439852 285776 442906 285832
rect 442962 285776 442967 285832
rect 439852 285774 442967 285776
rect 442901 285771 442967 285774
rect 583520 285276 584960 285516
rect 57329 283114 57395 283117
rect 440601 283114 440667 283117
rect 57329 283112 60076 283114
rect 57329 283056 57334 283112
rect 57390 283056 60076 283112
rect 57329 283054 60076 283056
rect 439852 283112 440667 283114
rect 439852 283056 440606 283112
rect 440662 283056 440667 283112
rect 439852 283054 440667 283056
rect 57329 283051 57395 283054
rect 440601 283051 440667 283054
rect 55857 280394 55923 280397
rect 55857 280392 60076 280394
rect 55857 280336 55862 280392
rect 55918 280336 60076 280392
rect 55857 280334 60076 280336
rect 55857 280331 55923 280334
rect -960 279972 480 280212
rect 442809 279714 442875 279717
rect 439852 279712 442875 279714
rect 439852 279656 442814 279712
rect 442870 279656 442875 279712
rect 439852 279654 442875 279656
rect 442809 279651 442875 279654
rect 57329 277674 57395 277677
rect 57329 277672 60076 277674
rect 57329 277616 57334 277672
rect 57390 277616 60076 277672
rect 57329 277614 60076 277616
rect 57329 277611 57395 277614
rect 442533 276994 442599 276997
rect 439852 276992 442599 276994
rect 439852 276936 442538 276992
rect 442594 276936 442599 276992
rect 439852 276934 442599 276936
rect 442533 276931 442599 276934
rect 60590 274484 60596 274548
rect 60660 274484 60666 274548
rect 60598 274244 60658 274484
rect 442901 274274 442967 274277
rect 439852 274272 442967 274274
rect 439852 274216 442906 274272
rect 442962 274216 442967 274272
rect 439852 274214 442967 274216
rect 442901 274211 442967 274214
rect 580717 272234 580783 272237
rect 583520 272234 584960 272324
rect 580717 272232 584960 272234
rect 580717 272176 580722 272232
rect 580778 272176 584960 272232
rect 580717 272174 584960 272176
rect 580717 272171 580783 272174
rect 583520 272084 584960 272174
rect 57329 271554 57395 271557
rect 442901 271554 442967 271557
rect 57329 271552 60076 271554
rect 57329 271496 57334 271552
rect 57390 271496 60076 271552
rect 57329 271494 60076 271496
rect 439852 271552 442967 271554
rect 439852 271496 442906 271552
rect 442962 271496 442967 271552
rect 439852 271494 442967 271496
rect 57329 271491 57395 271494
rect 442901 271491 442967 271494
rect 56593 268834 56659 268837
rect 56593 268832 60076 268834
rect 56593 268776 56598 268832
rect 56654 268776 60076 268832
rect 56593 268774 60076 268776
rect 56593 268771 56659 268774
rect 442901 268154 442967 268157
rect 439852 268152 442967 268154
rect 439852 268096 442906 268152
rect 442962 268096 442967 268152
rect 439852 268094 442967 268096
rect 442901 268091 442967 268094
rect -960 267202 480 267292
rect 3877 267202 3943 267205
rect -960 267200 3943 267202
rect -960 267144 3882 267200
rect 3938 267144 3943 267200
rect -960 267142 3943 267144
rect -960 267052 480 267142
rect 3877 267139 3943 267142
rect 57421 266114 57487 266117
rect 57421 266112 60076 266114
rect 57421 266056 57426 266112
rect 57482 266056 60076 266112
rect 57421 266054 60076 266056
rect 57421 266051 57487 266054
rect 442901 265434 442967 265437
rect 439852 265432 442967 265434
rect 439852 265376 442906 265432
rect 442962 265376 442967 265432
rect 439852 265374 442967 265376
rect 442901 265371 442967 265374
rect 57421 262714 57487 262717
rect 442901 262714 442967 262717
rect 57421 262712 60076 262714
rect 57421 262656 57426 262712
rect 57482 262656 60076 262712
rect 57421 262654 60076 262656
rect 439852 262712 442967 262714
rect 439852 262656 442906 262712
rect 442962 262656 442967 262712
rect 439852 262654 442967 262656
rect 57421 262651 57487 262654
rect 442901 262651 442967 262654
rect 57329 259994 57395 259997
rect 57329 259992 60076 259994
rect 57329 259936 57334 259992
rect 57390 259936 60076 259992
rect 57329 259934 60076 259936
rect 57329 259931 57395 259934
rect 442901 259314 442967 259317
rect 439852 259312 442967 259314
rect 439852 259256 442906 259312
rect 442962 259256 442967 259312
rect 439852 259254 442967 259256
rect 442901 259251 442967 259254
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect 58617 257274 58683 257277
rect 58617 257272 60076 257274
rect 58617 257216 58622 257272
rect 58678 257216 60076 257272
rect 58617 257214 60076 257216
rect 58617 257211 58683 257214
rect 442533 256594 442599 256597
rect 439852 256592 442599 256594
rect 439852 256536 442538 256592
rect 442594 256536 442599 256592
rect 439852 256534 442599 256536
rect 442533 256531 442599 256534
rect 57421 254554 57487 254557
rect 57421 254552 60076 254554
rect 57421 254496 57426 254552
rect 57482 254496 60076 254552
rect 57421 254494 60076 254496
rect 57421 254491 57487 254494
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 442349 253874 442415 253877
rect 439852 253872 442415 253874
rect 439852 253816 442354 253872
rect 442410 253816 442415 253872
rect 439852 253814 442415 253816
rect 442349 253811 442415 253814
rect 56869 251154 56935 251157
rect 442901 251154 442967 251157
rect 56869 251152 60076 251154
rect 56869 251096 56874 251152
rect 56930 251096 60076 251152
rect 56869 251094 60076 251096
rect 439852 251152 442967 251154
rect 439852 251096 442906 251152
rect 442962 251096 442967 251152
rect 439852 251094 442967 251096
rect 56869 251091 56935 251094
rect 442901 251091 442967 251094
rect 57421 248434 57487 248437
rect 57421 248432 60076 248434
rect 57421 248376 57426 248432
rect 57482 248376 60076 248432
rect 57421 248374 60076 248376
rect 57421 248371 57487 248374
rect 442717 247754 442783 247757
rect 439852 247752 442783 247754
rect 439852 247696 442722 247752
rect 442778 247696 442783 247752
rect 439852 247694 442783 247696
rect 442717 247691 442783 247694
rect 58525 245714 58591 245717
rect 58525 245712 60076 245714
rect 58525 245656 58530 245712
rect 58586 245656 60076 245712
rect 58525 245654 60076 245656
rect 58525 245651 58591 245654
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 442901 245034 442967 245037
rect 439852 245032 442967 245034
rect 439852 244976 442906 245032
rect 442962 244976 442967 245032
rect 439852 244974 442967 244976
rect 442901 244971 442967 244974
rect 57329 242994 57395 242997
rect 57329 242992 60076 242994
rect 57329 242936 57334 242992
rect 57390 242936 60076 242992
rect 57329 242934 60076 242936
rect 57329 242931 57395 242934
rect 440601 242314 440667 242317
rect 439852 242312 440667 242314
rect 439852 242256 440606 242312
rect 440662 242256 440667 242312
rect 439852 242254 440667 242256
rect 440601 242251 440667 242254
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 57329 239594 57395 239597
rect 442717 239594 442783 239597
rect 57329 239592 60076 239594
rect 57329 239536 57334 239592
rect 57390 239536 60076 239592
rect 57329 239534 60076 239536
rect 439852 239592 442783 239594
rect 439852 239536 442722 239592
rect 442778 239536 442783 239592
rect 439852 239534 442783 239536
rect 57329 239531 57395 239534
rect 442717 239531 442783 239534
rect 57881 236874 57947 236877
rect 57881 236872 60076 236874
rect 57881 236816 57886 236872
rect 57942 236816 60076 236872
rect 57881 236814 60076 236816
rect 57881 236811 57947 236814
rect 442901 236194 442967 236197
rect 439852 236192 442967 236194
rect 439852 236136 442906 236192
rect 442962 236136 442967 236192
rect 439852 236134 442967 236136
rect 442901 236131 442967 236134
rect 57237 234154 57303 234157
rect 57237 234152 60076 234154
rect 57237 234096 57242 234152
rect 57298 234096 60076 234152
rect 57237 234094 60076 234096
rect 57237 234091 57303 234094
rect 442901 233474 442967 233477
rect 439852 233472 442967 233474
rect 439852 233416 442906 233472
rect 442962 233416 442967 233472
rect 439852 233414 442967 233416
rect 442901 233411 442967 233414
rect 583520 232386 584960 232476
rect 583342 232326 584960 232386
rect 583342 232250 583402 232326
rect 583520 232250 584960 232326
rect 583342 232236 584960 232250
rect 583342 232190 583586 232236
rect 450486 231916 450492 231980
rect 450556 231978 450562 231980
rect 583526 231978 583586 232190
rect 450556 231918 583586 231978
rect 450556 231916 450562 231918
rect 57329 230754 57395 230757
rect 442901 230754 442967 230757
rect 57329 230752 60076 230754
rect 57329 230696 57334 230752
rect 57390 230696 60076 230752
rect 57329 230694 60076 230696
rect 439852 230752 442967 230754
rect 439852 230696 442906 230752
rect 442962 230696 442967 230752
rect 439852 230694 442967 230696
rect 57329 230691 57395 230694
rect 442901 230691 442967 230694
rect -960 227884 480 228124
rect 57881 228034 57947 228037
rect 57881 228032 60076 228034
rect 57881 227976 57886 228032
rect 57942 227976 60076 228032
rect 57881 227974 60076 227976
rect 57881 227971 57947 227974
rect 442901 227354 442967 227357
rect 439852 227352 442967 227354
rect 439852 227296 442906 227352
rect 442962 227296 442967 227352
rect 439852 227294 442967 227296
rect 442901 227291 442967 227294
rect 57881 225314 57947 225317
rect 57881 225312 60076 225314
rect 57881 225256 57886 225312
rect 57942 225256 60076 225312
rect 57881 225254 60076 225256
rect 57881 225251 57947 225254
rect 441061 224634 441127 224637
rect 439852 224632 441127 224634
rect 439852 224576 441066 224632
rect 441122 224576 441127 224632
rect 439852 224574 441127 224576
rect 441061 224571 441127 224574
rect 57881 222594 57947 222597
rect 57881 222592 60076 222594
rect 57881 222536 57886 222592
rect 57942 222536 60076 222592
rect 57881 222534 60076 222536
rect 57881 222531 57947 222534
rect 442625 221914 442691 221917
rect 439852 221912 442691 221914
rect 439852 221856 442630 221912
rect 442686 221856 442691 221912
rect 439852 221854 442691 221856
rect 442625 221851 442691 221854
rect 57881 219194 57947 219197
rect 442901 219194 442967 219197
rect 57881 219192 60076 219194
rect 57881 219136 57886 219192
rect 57942 219136 60076 219192
rect 57881 219134 60076 219136
rect 439852 219192 442967 219194
rect 439852 219136 442906 219192
rect 442962 219136 442967 219192
rect 439852 219134 442967 219136
rect 57881 219131 57947 219134
rect 442901 219131 442967 219134
rect 579981 219058 580047 219061
rect 583520 219058 584960 219148
rect 579981 219056 584960 219058
rect 579981 219000 579986 219056
rect 580042 219000 584960 219056
rect 579981 218998 584960 219000
rect 579981 218995 580047 218998
rect 583520 218908 584960 218998
rect 56593 216474 56659 216477
rect 56593 216472 60076 216474
rect 56593 216416 56598 216472
rect 56654 216416 60076 216472
rect 56593 216414 60076 216416
rect 56593 216411 56659 216414
rect 442901 215794 442967 215797
rect 439852 215792 442967 215794
rect 439852 215736 442906 215792
rect 442962 215736 442967 215792
rect 439852 215734 442967 215736
rect 442901 215731 442967 215734
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 60598 213212 60658 213724
rect 60590 213148 60596 213212
rect 60660 213148 60666 213212
rect 442717 213074 442783 213077
rect 439852 213072 442783 213074
rect 439852 213016 442722 213072
rect 442778 213016 442783 213072
rect 439852 213014 442783 213016
rect 442717 213011 442783 213014
rect 57881 211034 57947 211037
rect 57881 211032 60076 211034
rect 57881 210976 57886 211032
rect 57942 210976 60076 211032
rect 57881 210974 60076 210976
rect 57881 210971 57947 210974
rect 442717 210354 442783 210357
rect 439852 210352 442783 210354
rect 439852 210296 442722 210352
rect 442778 210296 442783 210352
rect 439852 210294 442783 210296
rect 442717 210291 442783 210294
rect 57697 207634 57763 207637
rect 442441 207634 442507 207637
rect 57697 207632 60076 207634
rect 57697 207576 57702 207632
rect 57758 207576 60076 207632
rect 57697 207574 60076 207576
rect 439852 207632 442507 207634
rect 439852 207576 442446 207632
rect 442502 207576 442507 207632
rect 439852 207574 442507 207576
rect 57697 207571 57763 207574
rect 442441 207571 442507 207574
rect 580809 205730 580875 205733
rect 583520 205730 584960 205820
rect 580809 205728 584960 205730
rect 580809 205672 580814 205728
rect 580870 205672 584960 205728
rect 580809 205670 584960 205672
rect 580809 205667 580875 205670
rect 583520 205580 584960 205670
rect 57697 204914 57763 204917
rect 57697 204912 60076 204914
rect 57697 204856 57702 204912
rect 57758 204856 60076 204912
rect 57697 204854 60076 204856
rect 57697 204851 57763 204854
rect 442901 204234 442967 204237
rect 439852 204232 442967 204234
rect 439852 204176 442906 204232
rect 442962 204176 442967 204232
rect 439852 204174 442967 204176
rect 442901 204171 442967 204174
rect 3141 202874 3207 202877
rect 36486 202874 36492 202876
rect 3141 202872 36492 202874
rect 3141 202816 3146 202872
rect 3202 202816 36492 202872
rect 3141 202814 36492 202816
rect 3141 202811 3207 202814
rect 36486 202812 36492 202814
rect 36556 202812 36562 202876
rect 57881 202194 57947 202197
rect 57881 202192 60076 202194
rect 57881 202136 57886 202192
rect 57942 202136 60076 202192
rect 57881 202134 60076 202136
rect 57881 202131 57947 202134
rect -960 201922 480 202012
rect 3141 201922 3207 201925
rect -960 201920 3207 201922
rect -960 201864 3146 201920
rect 3202 201864 3207 201920
rect -960 201862 3207 201864
rect -960 201772 480 201862
rect 3141 201859 3207 201862
rect 442901 201514 442967 201517
rect 439852 201512 442967 201514
rect 439852 201456 442906 201512
rect 442962 201456 442967 201512
rect 439852 201454 442967 201456
rect 442901 201451 442967 201454
rect 56593 198794 56659 198797
rect 442901 198794 442967 198797
rect 56593 198792 60076 198794
rect 56593 198736 56598 198792
rect 56654 198736 60076 198792
rect 56593 198734 60076 198736
rect 439852 198792 442967 198794
rect 439852 198736 442906 198792
rect 442962 198736 442967 198792
rect 439852 198734 442967 198736
rect 56593 198731 56659 198734
rect 442901 198731 442967 198734
rect 57697 196074 57763 196077
rect 57697 196072 60076 196074
rect 57697 196016 57702 196072
rect 57758 196016 60076 196072
rect 57697 196014 60076 196016
rect 57697 196011 57763 196014
rect 442901 195394 442967 195397
rect 439852 195392 442967 195394
rect 439852 195336 442906 195392
rect 442962 195336 442967 195392
rect 439852 195334 442967 195336
rect 442901 195331 442967 195334
rect 57697 193354 57763 193357
rect 57697 193352 60076 193354
rect 57697 193296 57702 193352
rect 57758 193296 60076 193352
rect 57697 193294 60076 193296
rect 57697 193291 57763 193294
rect 442901 192674 442967 192677
rect 439852 192672 442967 192674
rect 439852 192616 442906 192672
rect 442962 192616 442967 192672
rect 439852 192614 442967 192616
rect 442901 192611 442967 192614
rect 580717 192538 580783 192541
rect 583520 192538 584960 192628
rect 580717 192536 584960 192538
rect 580717 192480 580722 192536
rect 580778 192480 584960 192536
rect 580717 192478 584960 192480
rect 580717 192475 580783 192478
rect 583520 192388 584960 192478
rect 56869 190634 56935 190637
rect 56869 190632 60076 190634
rect 56869 190576 56874 190632
rect 56930 190576 60076 190632
rect 56869 190574 60076 190576
rect 56869 190571 56935 190574
rect 441153 189954 441219 189957
rect 439852 189952 441219 189954
rect 439852 189896 441158 189952
rect 441214 189896 441219 189952
rect 439852 189894 441219 189896
rect 441153 189891 441219 189894
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 57697 187234 57763 187237
rect 442625 187234 442691 187237
rect 57697 187232 60076 187234
rect 57697 187176 57702 187232
rect 57758 187176 60076 187232
rect 57697 187174 60076 187176
rect 439852 187232 442691 187234
rect 439852 187176 442630 187232
rect 442686 187176 442691 187232
rect 439852 187174 442691 187176
rect 57697 187171 57763 187174
rect 442625 187171 442691 187174
rect 57697 184514 57763 184517
rect 57697 184512 60076 184514
rect 57697 184456 57702 184512
rect 57758 184456 60076 184512
rect 57697 184454 60076 184456
rect 57697 184451 57763 184454
rect 441245 183834 441311 183837
rect 439852 183832 441311 183834
rect 439852 183776 441250 183832
rect 441306 183776 441311 183832
rect 439852 183774 441311 183776
rect 441245 183771 441311 183774
rect 57697 181794 57763 181797
rect 57697 181792 60076 181794
rect 57697 181736 57702 181792
rect 57758 181736 60076 181792
rect 57697 181734 60076 181736
rect 57697 181731 57763 181734
rect 442901 181114 442967 181117
rect 439852 181112 442967 181114
rect 439852 181056 442906 181112
rect 442962 181056 442967 181112
rect 439852 181054 442967 181056
rect 442901 181051 442967 181054
rect 60590 179284 60596 179348
rect 60660 179284 60666 179348
rect 60598 179044 60658 179284
rect 580901 179210 580967 179213
rect 583520 179210 584960 179300
rect 580901 179208 584960 179210
rect 580901 179152 580906 179208
rect 580962 179152 584960 179208
rect 580901 179150 584960 179152
rect 580901 179147 580967 179150
rect 583520 179060 584960 179150
rect 442901 178394 442967 178397
rect 439852 178392 442967 178394
rect 439852 178336 442906 178392
rect 442962 178336 442967 178392
rect 439852 178334 442967 178336
rect 442901 178331 442967 178334
rect -960 175796 480 176036
rect 57881 175674 57947 175677
rect 442717 175674 442783 175677
rect 57881 175672 60076 175674
rect 57881 175616 57886 175672
rect 57942 175616 60076 175672
rect 57881 175614 60076 175616
rect 439852 175672 442783 175674
rect 439852 175616 442722 175672
rect 442778 175616 442783 175672
rect 439852 175614 442783 175616
rect 57881 175611 57947 175614
rect 442717 175611 442783 175614
rect 57697 172954 57763 172957
rect 57697 172952 60076 172954
rect 57697 172896 57702 172952
rect 57758 172896 60076 172952
rect 57697 172894 60076 172896
rect 57697 172891 57763 172894
rect 442901 172274 442967 172277
rect 439852 172272 442967 172274
rect 439852 172216 442906 172272
rect 442962 172216 442967 172272
rect 439852 172214 442967 172216
rect 442901 172211 442967 172214
rect 57881 170234 57947 170237
rect 57881 170232 60076 170234
rect 57881 170176 57886 170232
rect 57942 170176 60076 170232
rect 57881 170174 60076 170176
rect 57881 170171 57947 170174
rect 442901 169554 442967 169557
rect 439852 169552 442967 169554
rect 439852 169496 442906 169552
rect 442962 169496 442967 169552
rect 439852 169494 442967 169496
rect 442901 169491 442967 169494
rect 57881 166834 57947 166837
rect 57881 166832 60076 166834
rect 57881 166776 57886 166832
rect 57942 166776 60076 166832
rect 57881 166774 60076 166776
rect 57881 166771 57947 166774
rect 439822 166290 439882 166804
rect 439957 166290 440023 166293
rect 439822 166288 440023 166290
rect 439822 166232 439962 166288
rect 440018 166232 440023 166288
rect 439822 166230 440023 166232
rect 439957 166227 440023 166230
rect 580625 165882 580691 165885
rect 583520 165882 584960 165972
rect 580625 165880 584960 165882
rect 580625 165824 580630 165880
rect 580686 165824 584960 165880
rect 580625 165822 584960 165824
rect 580625 165819 580691 165822
rect 583520 165732 584960 165822
rect 57881 164114 57947 164117
rect 442533 164114 442599 164117
rect 57881 164112 60076 164114
rect 57881 164056 57886 164112
rect 57942 164056 60076 164112
rect 57881 164054 60076 164056
rect 439852 164112 442599 164114
rect 439852 164056 442538 164112
rect 442594 164056 442599 164112
rect 439852 164054 442599 164056
rect 57881 164051 57947 164054
rect 442533 164051 442599 164054
rect -960 162890 480 162980
rect 3877 162890 3943 162893
rect -960 162888 3943 162890
rect -960 162832 3882 162888
rect 3938 162832 3943 162888
rect -960 162830 3943 162832
rect -960 162740 480 162830
rect 3877 162827 3943 162830
rect 60598 160852 60658 161364
rect 60590 160788 60596 160852
rect 60660 160788 60666 160852
rect 442901 160714 442967 160717
rect 439852 160712 442967 160714
rect 439852 160656 442906 160712
rect 442962 160656 442967 160712
rect 439852 160654 442967 160656
rect 442901 160651 442967 160654
rect 57145 158674 57211 158677
rect 57145 158672 60076 158674
rect 57145 158616 57150 158672
rect 57206 158616 60076 158672
rect 57145 158614 60076 158616
rect 57145 158611 57211 158614
rect 442717 157994 442783 157997
rect 439852 157992 442783 157994
rect 439852 157936 442722 157992
rect 442778 157936 442783 157992
rect 439852 157934 442783 157936
rect 442717 157931 442783 157934
rect 57881 155274 57947 155277
rect 442625 155274 442691 155277
rect 57881 155272 60076 155274
rect 57881 155216 57886 155272
rect 57942 155216 60076 155272
rect 57881 155214 60076 155216
rect 439852 155272 442691 155274
rect 439852 155216 442630 155272
rect 442686 155216 442691 155272
rect 439852 155214 442691 155216
rect 57881 155211 57947 155214
rect 442625 155211 442691 155214
rect 580533 152690 580599 152693
rect 583520 152690 584960 152780
rect 580533 152688 584960 152690
rect 580533 152632 580538 152688
rect 580594 152632 584960 152688
rect 580533 152630 584960 152632
rect 580533 152627 580599 152630
rect 57881 152554 57947 152557
rect 57881 152552 60076 152554
rect 57881 152496 57886 152552
rect 57942 152496 60076 152552
rect 583520 152540 584960 152630
rect 57881 152494 60076 152496
rect 57881 152491 57947 152494
rect 439497 152418 439563 152421
rect 439454 152416 439563 152418
rect 439454 152360 439502 152416
rect 439558 152360 439563 152416
rect 439454 152355 439563 152360
rect 439454 151844 439514 152355
rect -960 149834 480 149924
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 57881 149834 57947 149837
rect 57881 149832 60076 149834
rect 57881 149776 57886 149832
rect 57942 149776 60076 149832
rect 57881 149774 60076 149776
rect 57881 149771 57947 149774
rect 442901 149154 442967 149157
rect 439852 149152 442967 149154
rect 439852 149096 442906 149152
rect 442962 149096 442967 149152
rect 439852 149094 442967 149096
rect 442901 149091 442967 149094
rect 57881 147114 57947 147117
rect 57881 147112 60076 147114
rect 57881 147056 57886 147112
rect 57942 147056 60076 147112
rect 57881 147054 60076 147056
rect 57881 147051 57947 147054
rect 442809 146434 442875 146437
rect 439852 146432 442875 146434
rect 439852 146376 442814 146432
rect 442870 146376 442875 146432
rect 439852 146374 442875 146376
rect 442809 146371 442875 146374
rect 57053 143714 57119 143717
rect 442901 143714 442967 143717
rect 57053 143712 60076 143714
rect 57053 143656 57058 143712
rect 57114 143656 60076 143712
rect 57053 143654 60076 143656
rect 439852 143712 442967 143714
rect 439852 143656 442906 143712
rect 442962 143656 442967 143712
rect 439852 143654 442967 143656
rect 57053 143651 57119 143654
rect 442901 143651 442967 143654
rect 57881 140994 57947 140997
rect 57881 140992 60076 140994
rect 57881 140936 57886 140992
rect 57942 140936 60076 140992
rect 57881 140934 60076 140936
rect 57881 140931 57947 140934
rect 442901 140314 442967 140317
rect 439852 140312 442967 140314
rect 439852 140256 442906 140312
rect 442962 140256 442967 140312
rect 439852 140254 442967 140256
rect 442901 140251 442967 140254
rect 583520 139362 584960 139452
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 59261 138274 59327 138277
rect 59261 138272 60076 138274
rect 59261 138216 59266 138272
rect 59322 138216 60076 138272
rect 59261 138214 60076 138216
rect 59261 138211 59327 138214
rect 453246 138076 453252 138140
rect 453316 138138 453322 138140
rect 583526 138138 583586 139166
rect 453316 138078 583586 138138
rect 453316 138076 453322 138078
rect 442717 137594 442783 137597
rect 439852 137592 442783 137594
rect 439852 137536 442722 137592
rect 442778 137536 442783 137592
rect 439852 137534 442783 137536
rect 442717 137531 442783 137534
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 57881 135554 57947 135557
rect 57881 135552 60076 135554
rect 57881 135496 57886 135552
rect 57942 135496 60076 135552
rect 57881 135494 60076 135496
rect 57881 135491 57947 135494
rect 442901 134874 442967 134877
rect 439852 134872 442967 134874
rect 439852 134816 442906 134872
rect 442962 134816 442967 134872
rect 439852 134814 442967 134816
rect 442901 134811 442967 134814
rect 57881 132154 57947 132157
rect 442901 132154 442967 132157
rect 57881 132152 60076 132154
rect 57881 132096 57886 132152
rect 57942 132096 60076 132152
rect 57881 132094 60076 132096
rect 439852 132152 442967 132154
rect 439852 132096 442906 132152
rect 442962 132096 442967 132152
rect 439852 132094 442967 132096
rect 57881 132091 57947 132094
rect 442901 132091 442967 132094
rect 57881 129434 57947 129437
rect 57881 129432 60076 129434
rect 57881 129376 57886 129432
rect 57942 129376 60076 129432
rect 57881 129374 60076 129376
rect 57881 129371 57947 129374
rect 442901 128754 442967 128757
rect 439852 128752 442967 128754
rect 439852 128696 442906 128752
rect 442962 128696 442967 128752
rect 439852 128694 442967 128696
rect 442901 128691 442967 128694
rect 56961 126714 57027 126717
rect 56961 126712 60076 126714
rect 56961 126656 56966 126712
rect 57022 126656 60076 126712
rect 56961 126654 60076 126656
rect 56961 126651 57027 126654
rect 583520 126034 584960 126124
rect 439822 125762 439882 126004
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 441521 125762 441587 125765
rect 439822 125760 441587 125762
rect 439822 125704 441526 125760
rect 441582 125704 441587 125760
rect 439822 125702 441587 125704
rect 441521 125699 441587 125702
rect 468334 125564 468340 125628
rect 468404 125626 468410 125628
rect 583526 125626 583586 125838
rect 468404 125566 583586 125626
rect 468404 125564 468410 125566
rect -960 123572 480 123812
rect 57881 123314 57947 123317
rect 57881 123312 60076 123314
rect 57881 123256 57886 123312
rect 57942 123256 60076 123312
rect 57881 123254 60076 123256
rect 57881 123251 57947 123254
rect 439822 122906 439882 123284
rect 441521 122906 441587 122909
rect 439822 122904 441587 122906
rect 439822 122848 441526 122904
rect 441582 122848 441587 122904
rect 439822 122846 441587 122848
rect 441521 122843 441587 122846
rect 57881 120594 57947 120597
rect 57881 120592 60076 120594
rect 57881 120536 57886 120592
rect 57942 120536 60076 120592
rect 57881 120534 60076 120536
rect 57881 120531 57947 120534
rect 439822 119370 439882 119884
rect 441521 119370 441587 119373
rect 439822 119368 441587 119370
rect 439822 119312 441526 119368
rect 441582 119312 441587 119368
rect 439822 119310 441587 119312
rect 441521 119307 441587 119310
rect 57881 117874 57947 117877
rect 57881 117872 60076 117874
rect 57881 117816 57886 117872
rect 57942 117816 60076 117872
rect 57881 117814 60076 117816
rect 57881 117811 57947 117814
rect 439822 116650 439882 117164
rect 441521 116650 441587 116653
rect 439822 116648 441587 116650
rect 439822 116592 441526 116648
rect 441582 116592 441587 116648
rect 439822 116590 441587 116592
rect 441521 116587 441587 116590
rect 57881 115154 57947 115157
rect 57881 115152 60076 115154
rect 57881 115096 57886 115152
rect 57942 115096 60076 115152
rect 57881 115094 60076 115096
rect 57881 115091 57947 115094
rect 441521 114474 441587 114477
rect 439852 114472 441587 114474
rect 439852 114416 441526 114472
rect 441582 114416 441587 114472
rect 439852 114414 441587 114416
rect 441521 114411 441587 114414
rect 579981 112842 580047 112845
rect 583520 112842 584960 112932
rect 579981 112840 584960 112842
rect 579981 112784 579986 112840
rect 580042 112784 584960 112840
rect 579981 112782 584960 112784
rect 579981 112779 580047 112782
rect 583520 112692 584960 112782
rect 3141 111754 3207 111757
rect 32254 111754 32260 111756
rect 3141 111752 32260 111754
rect 3141 111696 3146 111752
rect 3202 111696 32260 111752
rect 3141 111694 32260 111696
rect 3141 111691 3207 111694
rect 32254 111692 32260 111694
rect 32324 111692 32330 111756
rect 59721 111754 59787 111757
rect 59721 111752 60076 111754
rect 59721 111696 59726 111752
rect 59782 111696 60076 111752
rect 59721 111694 60076 111696
rect 59721 111691 59787 111694
rect 439822 111210 439882 111724
rect 441521 111210 441587 111213
rect 439822 111208 441587 111210
rect 439822 111152 441526 111208
rect 441582 111152 441587 111208
rect 439822 111150 441587 111152
rect 441521 111147 441587 111150
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 59261 109034 59327 109037
rect 59261 109032 60076 109034
rect 59261 108976 59266 109032
rect 59322 108976 60076 109032
rect 59261 108974 60076 108976
rect 59261 108971 59327 108974
rect 439822 107810 439882 108324
rect 441521 107810 441587 107813
rect 439822 107808 441587 107810
rect 439822 107752 441526 107808
rect 441582 107752 441587 107808
rect 439822 107750 441587 107752
rect 441521 107747 441587 107750
rect 57881 106314 57947 106317
rect 57881 106312 60076 106314
rect 57881 106256 57886 106312
rect 57942 106256 60076 106312
rect 57881 106254 60076 106256
rect 57881 106251 57947 106254
rect 439822 105090 439882 105604
rect 441521 105090 441587 105093
rect 439822 105088 441587 105090
rect 439822 105032 441526 105088
rect 441582 105032 441587 105088
rect 439822 105030 441587 105032
rect 441521 105027 441587 105030
rect 56593 103594 56659 103597
rect 56593 103592 60076 103594
rect 56593 103536 56598 103592
rect 56654 103536 60076 103592
rect 56593 103534 60076 103536
rect 56593 103531 56659 103534
rect 441521 103458 441587 103461
rect 439822 103456 441587 103458
rect 439822 103400 441526 103456
rect 441582 103400 441587 103456
rect 439822 103398 441587 103400
rect 439822 102884 439882 103398
rect 441521 103395 441587 103398
rect 57881 100194 57947 100197
rect 57881 100192 60076 100194
rect 57881 100136 57886 100192
rect 57942 100136 60076 100192
rect 57881 100134 60076 100136
rect 57881 100131 57947 100134
rect 439822 99650 439882 100164
rect 441521 99650 441587 99653
rect 439822 99648 441587 99650
rect 439822 99592 441526 99648
rect 441582 99592 441587 99648
rect 439822 99590 441587 99592
rect 441521 99587 441587 99590
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 22686 97882 22692 97884
rect 6870 97822 22692 97882
rect -960 97610 480 97700
rect 6870 97610 6930 97822
rect 22686 97820 22692 97822
rect 22756 97820 22762 97884
rect -960 97550 6930 97610
rect -960 97460 480 97550
rect 58433 97474 58499 97477
rect 58433 97472 60076 97474
rect 58433 97416 58438 97472
rect 58494 97416 60076 97472
rect 58433 97414 60076 97416
rect 58433 97411 58499 97414
rect 439822 96661 439882 96764
rect 439822 96656 439931 96661
rect 439822 96600 439870 96656
rect 439926 96600 439931 96656
rect 439822 96598 439931 96600
rect 439865 96595 439931 96598
rect 57881 94754 57947 94757
rect 57881 94752 60076 94754
rect 57881 94696 57886 94752
rect 57942 94696 60076 94752
rect 57881 94694 60076 94696
rect 57881 94691 57947 94694
rect 439822 93941 439882 94044
rect 439773 93936 439882 93941
rect 439773 93880 439778 93936
rect 439834 93880 439882 93936
rect 439773 93878 439882 93880
rect 439773 93875 439839 93878
rect 58341 91354 58407 91357
rect 58341 91352 60076 91354
rect 58341 91296 58346 91352
rect 58402 91296 60076 91352
rect 58341 91294 60076 91296
rect 58341 91291 58407 91294
rect 439822 91218 439882 91324
rect 441521 91218 441587 91221
rect 439822 91216 441587 91218
rect 439822 91160 441526 91216
rect 441582 91160 441587 91216
rect 439822 91158 441587 91160
rect 441521 91155 441587 91158
rect 57881 88634 57947 88637
rect 57881 88632 60076 88634
rect 57881 88576 57886 88632
rect 57942 88576 60076 88632
rect 57881 88574 60076 88576
rect 57881 88571 57947 88574
rect 439822 87410 439882 87924
rect 441521 87410 441587 87413
rect 439822 87408 441587 87410
rect 439822 87352 441526 87408
rect 441582 87352 441587 87408
rect 439822 87350 441587 87352
rect 441521 87347 441587 87350
rect 580533 86186 580599 86189
rect 583520 86186 584960 86276
rect 580533 86184 584960 86186
rect 580533 86128 580538 86184
rect 580594 86128 584960 86184
rect 580533 86126 584960 86128
rect 580533 86123 580599 86126
rect 583520 86036 584960 86126
rect 57881 85914 57947 85917
rect 57881 85912 60076 85914
rect 57881 85856 57886 85912
rect 57942 85856 60076 85912
rect 57881 85854 60076 85856
rect 57881 85851 57947 85854
rect 441337 85234 441403 85237
rect 439852 85232 441403 85234
rect 439852 85176 441342 85232
rect 441398 85176 441403 85232
rect 439852 85174 441403 85176
rect 441337 85171 441403 85174
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 58249 83194 58315 83197
rect 58249 83192 60076 83194
rect 58249 83136 58254 83192
rect 58310 83136 60076 83192
rect 58249 83134 60076 83136
rect 58249 83131 58315 83134
rect 439822 81970 439882 82484
rect 441521 81970 441587 81973
rect 439822 81968 441587 81970
rect 439822 81912 441526 81968
rect 441582 81912 441587 81968
rect 439822 81910 441587 81912
rect 441521 81907 441587 81910
rect 59813 79794 59879 79797
rect 441521 79794 441587 79797
rect 59813 79792 60076 79794
rect 59813 79736 59818 79792
rect 59874 79736 60076 79792
rect 59813 79734 60076 79736
rect 439852 79792 441587 79794
rect 439852 79736 441526 79792
rect 441582 79736 441587 79792
rect 439852 79734 441587 79736
rect 59813 79731 59879 79734
rect 441521 79731 441587 79734
rect 56869 77074 56935 77077
rect 56869 77072 60076 77074
rect 56869 77016 56874 77072
rect 56930 77016 60076 77072
rect 56869 77014 60076 77016
rect 56869 77011 56935 77014
rect 441521 76394 441587 76397
rect 439852 76392 441587 76394
rect 439852 76336 441526 76392
rect 441582 76336 441587 76392
rect 439852 76334 441587 76336
rect 441521 76331 441587 76334
rect 58157 74354 58223 74357
rect 58157 74352 60076 74354
rect 58157 74296 58162 74352
rect 58218 74296 60076 74352
rect 58157 74294 60076 74296
rect 58157 74291 58223 74294
rect 439454 73133 439514 73644
rect 439454 73128 439563 73133
rect 439454 73072 439502 73128
rect 439558 73072 439563 73128
rect 439454 73070 439563 73072
rect 439497 73067 439563 73070
rect 580625 72994 580691 72997
rect 583520 72994 584960 73084
rect 580625 72992 584960 72994
rect 580625 72936 580630 72992
rect 580686 72936 584960 72992
rect 580625 72934 584960 72936
rect 580625 72931 580691 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 56777 71634 56843 71637
rect 56777 71632 60076 71634
rect 56777 71576 56782 71632
rect 56838 71576 60076 71632
rect 56777 71574 60076 71576
rect 56777 71571 56843 71574
rect 441429 70954 441495 70957
rect 439852 70952 441495 70954
rect 439852 70896 441434 70952
rect 441490 70896 441495 70952
rect 439852 70894 441495 70896
rect 441429 70891 441495 70894
rect 58065 68234 58131 68237
rect 58065 68232 60076 68234
rect 58065 68176 58070 68232
rect 58126 68176 60076 68232
rect 58065 68174 60076 68176
rect 58065 68171 58131 68174
rect 439822 67690 439882 68204
rect 440049 67690 440115 67693
rect 439822 67688 440115 67690
rect 439822 67632 440054 67688
rect 440110 67632 440115 67688
rect 439822 67630 440115 67632
rect 440049 67627 440115 67630
rect 56869 65514 56935 65517
rect 56869 65512 60076 65514
rect 56869 65456 56874 65512
rect 56930 65456 60076 65512
rect 56869 65454 60076 65456
rect 56869 65451 56935 65454
rect 440141 64834 440207 64837
rect 439852 64832 440207 64834
rect 439852 64776 440146 64832
rect 440202 64776 440207 64832
rect 439852 64774 440207 64776
rect 440141 64771 440207 64774
rect 59813 62794 59879 62797
rect 59813 62792 60076 62794
rect 59813 62736 59818 62792
rect 59874 62736 60076 62792
rect 59813 62734 60076 62736
rect 59813 62731 59879 62734
rect 439822 61570 439882 62084
rect 441521 61570 441587 61573
rect 439822 61568 441587 61570
rect 439822 61512 441526 61568
rect 441582 61512 441587 61568
rect 439822 61510 441587 61512
rect 441521 61507 441587 61510
rect 53097 61434 53163 61437
rect 560293 61434 560359 61437
rect 53097 61432 560359 61434
rect 53097 61376 53102 61432
rect 53158 61376 560298 61432
rect 560354 61376 560359 61432
rect 53097 61374 560359 61376
rect 53097 61371 53163 61374
rect 560293 61371 560359 61374
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2957 58578 3023 58581
rect -960 58576 3023 58578
rect -960 58520 2962 58576
rect 3018 58520 3023 58576
rect -960 58518 3023 58520
rect -960 58428 480 58518
rect 2957 58515 3023 58518
rect 219198 57836 219204 57900
rect 219268 57898 219274 57900
rect 381353 57898 381419 57901
rect 219268 57896 381419 57898
rect 219268 57840 381358 57896
rect 381414 57840 381419 57896
rect 219268 57838 381419 57840
rect 219268 57836 219274 57838
rect 381353 57835 381419 57838
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 342161 40626 342227 40629
rect 367686 40626 367692 40628
rect 342161 40624 367692 40626
rect 342161 40568 342166 40624
rect 342222 40568 367692 40624
rect 342161 40566 367692 40568
rect 342161 40563 342227 40566
rect 367686 40564 367692 40566
rect 367756 40564 367762 40628
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 152406 26828 152412 26892
rect 152476 26890 152482 26892
rect 237373 26890 237439 26893
rect 152476 26888 237439 26890
rect 152476 26832 237378 26888
rect 237434 26832 237439 26888
rect 152476 26830 237439 26832
rect 152476 26828 152482 26830
rect 237373 26827 237439 26830
rect 144821 24170 144887 24173
rect 219934 24170 219940 24172
rect 144821 24168 219940 24170
rect 144821 24112 144826 24168
rect 144882 24112 219940 24168
rect 144821 24110 219940 24112
rect 144821 24107 144887 24110
rect 219934 24108 219940 24110
rect 220004 24108 220010 24172
rect 252461 24170 252527 24173
rect 388110 24170 388116 24172
rect 252461 24168 388116 24170
rect 252461 24112 252466 24168
rect 252522 24112 388116 24168
rect 252461 24110 388116 24112
rect 252461 24107 252527 24110
rect 388110 24108 388116 24110
rect 388180 24108 388186 24172
rect 162761 21450 162827 21453
rect 269614 21450 269620 21452
rect 162761 21448 269620 21450
rect 162761 21392 162766 21448
rect 162822 21392 269620 21448
rect 162761 21390 269620 21392
rect 162761 21387 162827 21390
rect 269614 21388 269620 21390
rect 269684 21388 269690 21452
rect 137921 21314 137987 21317
rect 161974 21314 161980 21316
rect 137921 21312 161980 21314
rect 137921 21256 137926 21312
rect 137982 21256 161980 21312
rect 137921 21254 161980 21256
rect 137921 21251 137987 21254
rect 161974 21252 161980 21254
rect 162044 21252 162050 21316
rect 251766 21252 251772 21316
rect 251836 21314 251842 21316
rect 385033 21314 385099 21317
rect 251836 21312 385099 21314
rect 251836 21256 385038 21312
rect 385094 21256 385099 21312
rect 251836 21254 385099 21256
rect 251836 21252 251842 21254
rect 385033 21251 385099 21254
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 217961 18730 218027 18733
rect 384982 18730 384988 18732
rect 217961 18728 384988 18730
rect 217961 18672 217966 18728
rect 218022 18672 384988 18728
rect 217961 18670 384988 18672
rect 217961 18667 218027 18670
rect 384982 18668 384988 18670
rect 385052 18668 385058 18732
rect 119838 18532 119844 18596
rect 119908 18594 119914 18596
rect 380893 18594 380959 18597
rect 119908 18592 380959 18594
rect 119908 18536 380898 18592
rect 380954 18536 380959 18592
rect 119908 18534 380959 18536
rect 119908 18532 119914 18534
rect 380893 18531 380959 18534
rect 155861 17506 155927 17509
rect 240358 17506 240364 17508
rect 155861 17504 240364 17506
rect 155861 17448 155866 17504
rect 155922 17448 240364 17504
rect 155861 17446 240364 17448
rect 155861 17443 155927 17446
rect 240358 17444 240364 17446
rect 240428 17444 240434 17508
rect 155718 17308 155724 17372
rect 155788 17370 155794 17372
rect 281533 17370 281599 17373
rect 155788 17368 281599 17370
rect 155788 17312 281538 17368
rect 281594 17312 281599 17368
rect 155788 17310 281599 17312
rect 155788 17308 155794 17310
rect 281533 17307 281599 17310
rect 125358 17172 125364 17236
rect 125428 17234 125434 17236
rect 322933 17234 322999 17237
rect 125428 17232 322999 17234
rect 125428 17176 322938 17232
rect 322994 17176 322999 17232
rect 125428 17174 322999 17176
rect 125428 17172 125434 17174
rect 322933 17171 322999 17174
rect 222694 15812 222700 15876
rect 222764 15874 222770 15876
rect 246389 15874 246455 15877
rect 222764 15872 246455 15874
rect 222764 15816 246394 15872
rect 246450 15816 246455 15872
rect 222764 15814 246455 15816
rect 222764 15812 222770 15814
rect 246389 15811 246455 15814
rect 296621 15874 296687 15877
rect 313222 15874 313228 15876
rect 296621 15872 313228 15874
rect 296621 15816 296626 15872
rect 296682 15816 313228 15872
rect 296621 15814 313228 15816
rect 296621 15811 296687 15814
rect 313222 15812 313228 15814
rect 313292 15812 313298 15876
rect 332501 15874 332567 15877
rect 353886 15874 353892 15876
rect 332501 15872 353892 15874
rect 332501 15816 332506 15872
rect 332562 15816 353892 15872
rect 332501 15814 353892 15816
rect 332501 15811 332567 15814
rect 353886 15812 353892 15814
rect 353956 15812 353962 15876
rect 231761 14650 231827 14653
rect 363454 14650 363460 14652
rect 231761 14648 363460 14650
rect 231761 14592 231766 14648
rect 231822 14592 363460 14648
rect 231761 14590 363460 14592
rect 231761 14587 231827 14590
rect 363454 14588 363460 14590
rect 363524 14588 363530 14652
rect 106774 14452 106780 14516
rect 106844 14514 106850 14516
rect 240501 14514 240567 14517
rect 106844 14512 240567 14514
rect 106844 14456 240506 14512
rect 240562 14456 240567 14512
rect 106844 14454 240567 14456
rect 106844 14452 106850 14454
rect 240501 14451 240567 14454
rect 208894 13092 208900 13156
rect 208964 13154 208970 13156
rect 363505 13154 363571 13157
rect 208964 13152 363571 13154
rect 208964 13096 363510 13152
rect 363566 13096 363571 13152
rect 208964 13094 363571 13096
rect 208964 13092 208970 13094
rect 363505 13091 363571 13094
rect 139301 13018 139367 13021
rect 400806 13018 400812 13020
rect 139301 13016 400812 13018
rect 139301 12960 139306 13016
rect 139362 12960 400812 13016
rect 139301 12958 400812 12960
rect 139301 12955 139367 12958
rect 400806 12956 400812 12958
rect 400876 12956 400882 13020
rect 216581 12066 216647 12069
rect 242014 12066 242020 12068
rect 216581 12064 242020 12066
rect 216581 12008 216586 12064
rect 216642 12008 242020 12064
rect 216581 12006 242020 12008
rect 216581 12003 216647 12006
rect 242014 12004 242020 12006
rect 242084 12004 242090 12068
rect 166206 11868 166212 11932
rect 166276 11930 166282 11932
rect 307845 11930 307911 11933
rect 166276 11928 307911 11930
rect 166276 11872 307850 11928
rect 307906 11872 307911 11928
rect 166276 11870 307911 11872
rect 166276 11868 166282 11870
rect 307845 11867 307911 11870
rect 205541 11794 205607 11797
rect 228214 11794 228220 11796
rect 205541 11792 228220 11794
rect 205541 11736 205546 11792
rect 205602 11736 228220 11792
rect 205541 11734 228220 11736
rect 205541 11731 205607 11734
rect 228214 11732 228220 11734
rect 228284 11732 228290 11796
rect 237966 11732 237972 11796
rect 238036 11794 238042 11796
rect 390645 11794 390711 11797
rect 238036 11792 390711 11794
rect 238036 11736 390650 11792
rect 390706 11736 390711 11792
rect 238036 11734 390711 11736
rect 238036 11732 238042 11734
rect 390645 11731 390711 11734
rect 145925 11658 145991 11661
rect 322054 11658 322060 11660
rect 145925 11656 322060 11658
rect 145925 11600 145930 11656
rect 145986 11600 322060 11656
rect 145925 11598 322060 11600
rect 145925 11595 145991 11598
rect 322054 11596 322060 11598
rect 322124 11596 322130 11660
rect 253473 10978 253539 10981
rect 255814 10978 255820 10980
rect 253473 10976 255820 10978
rect 253473 10920 253478 10976
rect 253534 10920 255820 10976
rect 253473 10918 255820 10920
rect 253473 10915 253539 10918
rect 255814 10916 255820 10918
rect 255884 10916 255890 10980
rect 280654 10372 280660 10436
rect 280724 10434 280730 10436
rect 293677 10434 293743 10437
rect 280724 10432 293743 10434
rect 280724 10376 293682 10432
rect 293738 10376 293743 10432
rect 280724 10374 293743 10376
rect 280724 10372 280730 10374
rect 293677 10371 293743 10374
rect 327574 10372 327580 10436
rect 327644 10434 327650 10436
rect 373993 10434 374059 10437
rect 327644 10432 374059 10434
rect 327644 10376 373998 10432
rect 374054 10376 374059 10432
rect 327644 10374 374059 10376
rect 327644 10372 327650 10374
rect 373993 10371 374059 10374
rect 246246 10236 246252 10300
rect 246316 10298 246322 10300
rect 351637 10298 351703 10301
rect 246316 10296 351703 10298
rect 246316 10240 351642 10296
rect 351698 10240 351703 10296
rect 246316 10238 351703 10240
rect 246316 10236 246322 10238
rect 351637 10235 351703 10238
rect 336273 9618 336339 9621
rect 341190 9618 341196 9620
rect 336273 9616 341196 9618
rect 336273 9560 336278 9616
rect 336334 9560 341196 9616
rect 336273 9558 341196 9560
rect 336273 9555 336339 9558
rect 341190 9556 341196 9558
rect 341260 9556 341266 9620
rect 371693 9074 371759 9077
rect 389766 9074 389772 9076
rect 371693 9072 389772 9074
rect 371693 9016 371698 9072
rect 371754 9016 389772 9072
rect 371693 9014 389772 9016
rect 371693 9011 371759 9014
rect 389766 9012 389772 9014
rect 389836 9012 389842 9076
rect 344553 8938 344619 8941
rect 382222 8938 382228 8940
rect 344553 8936 382228 8938
rect 344553 8880 344558 8936
rect 344614 8880 382228 8936
rect 344553 8878 382228 8880
rect 344553 8875 344619 8878
rect 382222 8876 382228 8878
rect 382292 8876 382298 8940
rect 137134 7652 137140 7716
rect 137204 7714 137210 7716
rect 154205 7714 154271 7717
rect 137204 7712 154271 7714
rect 137204 7656 154210 7712
rect 154266 7656 154271 7712
rect 137204 7654 154271 7656
rect 137204 7652 137210 7654
rect 154205 7651 154271 7654
rect 54753 7578 54819 7581
rect 563237 7578 563303 7581
rect 54753 7576 563303 7578
rect 54753 7520 54758 7576
rect 54814 7520 563242 7576
rect 563298 7520 563303 7576
rect 54753 7518 563303 7520
rect 54753 7515 54819 7518
rect 563237 7515 563303 7518
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 244089 5674 244155 5677
rect 250294 5674 250300 5676
rect 244089 5672 250300 5674
rect 244089 5616 244094 5672
rect 244150 5616 250300 5672
rect 244089 5614 250300 5616
rect 244089 5611 244155 5614
rect 250294 5612 250300 5614
rect 250364 5612 250370 5676
rect 261753 5674 261819 5677
rect 266854 5674 266860 5676
rect 261753 5672 266860 5674
rect 261753 5616 261758 5672
rect 261814 5616 266860 5672
rect 261753 5614 266860 5616
rect 261753 5611 261819 5614
rect 266854 5612 266860 5614
rect 266924 5612 266930 5676
rect 332685 5674 332751 5677
rect 335854 5674 335860 5676
rect 332685 5672 335860 5674
rect 332685 5616 332690 5672
rect 332746 5616 335860 5672
rect 332685 5614 335860 5616
rect 332685 5611 332751 5614
rect 335854 5612 335860 5614
rect 335924 5612 335930 5676
rect 193213 4178 193279 4181
rect 197854 4178 197860 4180
rect 193213 4176 197860 4178
rect 193213 4120 193218 4176
rect 193274 4120 197860 4176
rect 193213 4118 197860 4120
rect 193213 4115 193279 4118
rect 197854 4116 197860 4118
rect 197924 4116 197930 4180
rect 230974 4116 230980 4180
rect 231044 4178 231050 4180
rect 235809 4178 235875 4181
rect 231044 4176 235875 4178
rect 231044 4120 235814 4176
rect 235870 4120 235875 4176
rect 231044 4118 235875 4120
rect 231044 4116 231050 4118
rect 235809 4115 235875 4118
rect 271086 4116 271092 4180
rect 271156 4178 271162 4180
rect 276013 4178 276079 4181
rect 271156 4176 276079 4178
rect 271156 4120 276018 4176
rect 276074 4120 276079 4176
rect 271156 4118 276079 4120
rect 271156 4116 271162 4118
rect 276013 4115 276079 4118
rect 277894 4116 277900 4180
rect 277964 4178 277970 4180
rect 279509 4178 279575 4181
rect 277964 4176 279575 4178
rect 277964 4120 279514 4176
rect 279570 4120 279575 4176
rect 277964 4118 279575 4120
rect 277964 4116 277970 4118
rect 279509 4115 279575 4118
rect 331806 4116 331812 4180
rect 331876 4178 331882 4180
rect 333881 4178 333947 4181
rect 331876 4176 333947 4178
rect 331876 4120 333886 4176
rect 333942 4120 333947 4176
rect 331876 4118 333947 4120
rect 331876 4116 331882 4118
rect 333881 4115 333947 4118
rect 72918 3980 72924 4044
rect 72988 4042 72994 4044
rect 109309 4042 109375 4045
rect 72988 4040 109375 4042
rect 72988 3984 109314 4040
rect 109370 3984 109375 4040
rect 72988 3982 109375 3984
rect 72988 3980 72994 3982
rect 109309 3979 109375 3982
rect 117589 4042 117655 4045
rect 298134 4042 298140 4044
rect 117589 4040 298140 4042
rect 117589 3984 117594 4040
rect 117650 3984 298140 4040
rect 117589 3982 298140 3984
rect 117589 3979 117655 3982
rect 298134 3980 298140 3982
rect 298204 3980 298210 4044
rect 393497 4042 393563 4045
rect 393814 4042 393820 4044
rect 393497 4040 393820 4042
rect 393497 3984 393502 4040
rect 393558 3984 393820 4040
rect 393497 3982 393820 3984
rect 393497 3979 393563 3982
rect 393814 3980 393820 3982
rect 393884 3980 393890 4044
rect 64321 3906 64387 3909
rect 442533 3906 442599 3909
rect 64321 3904 442599 3906
rect 64321 3848 64326 3904
rect 64382 3848 442538 3904
rect 442594 3848 442599 3904
rect 64321 3846 442599 3848
rect 64321 3843 64387 3846
rect 442533 3843 442599 3846
rect 45461 3770 45527 3773
rect 442717 3770 442783 3773
rect 45461 3768 442783 3770
rect 45461 3712 45466 3768
rect 45522 3712 442722 3768
rect 442778 3712 442783 3768
rect 45461 3710 442783 3712
rect 45461 3707 45527 3710
rect 442717 3707 442783 3710
rect 40677 3634 40743 3637
rect 442901 3634 442967 3637
rect 40677 3632 442967 3634
rect 40677 3576 40682 3632
rect 40738 3576 442906 3632
rect 442962 3576 442967 3632
rect 40677 3574 442967 3576
rect 40677 3571 40743 3574
rect 442901 3571 442967 3574
rect 34789 3498 34855 3501
rect 442257 3498 442323 3501
rect 34789 3496 442323 3498
rect 34789 3440 34794 3496
rect 34850 3440 442262 3496
rect 442318 3440 442323 3496
rect 34789 3438 442323 3440
rect 34789 3435 34855 3438
rect 442257 3435 442323 3438
rect 23013 3362 23079 3365
rect 442809 3362 442875 3365
rect 23013 3360 442875 3362
rect 23013 3304 23018 3360
rect 23074 3304 442814 3360
rect 442870 3304 442875 3360
rect 23013 3302 442875 3304
rect 23013 3299 23079 3302
rect 442809 3299 442875 3302
rect 73797 3226 73863 3229
rect 252502 3226 252508 3228
rect 73797 3224 252508 3226
rect 73797 3168 73802 3224
rect 73858 3168 252508 3224
rect 73797 3166 252508 3168
rect 73797 3163 73863 3166
rect 252502 3164 252508 3166
rect 252572 3164 252578 3228
rect 278998 3164 279004 3228
rect 279068 3226 279074 3228
rect 472249 3226 472315 3229
rect 279068 3224 472315 3226
rect 279068 3168 472254 3224
rect 472310 3168 472315 3224
rect 279068 3166 472315 3168
rect 279068 3164 279074 3166
rect 472249 3163 472315 3166
rect 57237 3090 57303 3093
rect 71681 3090 71747 3093
rect 57237 3088 71747 3090
rect 57237 3032 57242 3088
rect 57298 3032 71686 3088
rect 71742 3032 71747 3088
rect 57237 3030 71747 3032
rect 57237 3027 57303 3030
rect 71681 3027 71747 3030
rect 75678 3028 75684 3092
rect 75748 3090 75754 3092
rect 108113 3090 108179 3093
rect 118785 3090 118851 3093
rect 283782 3090 283788 3092
rect 75748 3088 108179 3090
rect 75748 3032 108118 3088
rect 108174 3032 108179 3088
rect 75748 3030 108179 3032
rect 75748 3028 75754 3030
rect 108113 3027 108179 3030
rect 108254 3030 118066 3090
rect 106917 2954 106983 2957
rect 108254 2954 108314 3030
rect 106917 2952 108314 2954
rect 106917 2896 106922 2952
rect 106978 2896 108314 2952
rect 106917 2894 108314 2896
rect 110505 2954 110571 2957
rect 118006 2954 118066 3030
rect 118785 3088 283788 3090
rect 118785 3032 118790 3088
rect 118846 3032 283788 3088
rect 118785 3030 283788 3032
rect 118785 3027 118851 3030
rect 283782 3028 283788 3030
rect 283852 3028 283858 3092
rect 304942 3028 304948 3092
rect 305012 3090 305018 3092
rect 305545 3090 305611 3093
rect 305012 3088 305611 3090
rect 305012 3032 305550 3088
rect 305606 3032 305611 3088
rect 305012 3030 305611 3032
rect 305012 3028 305018 3030
rect 305545 3027 305611 3030
rect 329833 3090 329899 3093
rect 330334 3090 330340 3092
rect 329833 3088 330340 3090
rect 329833 3032 329838 3088
rect 329894 3032 330340 3088
rect 329833 3030 330340 3032
rect 329833 3027 329899 3030
rect 330334 3028 330340 3030
rect 330404 3028 330410 3092
rect 350390 3028 350396 3092
rect 350460 3090 350466 3092
rect 583385 3090 583451 3093
rect 350460 3088 583451 3090
rect 350460 3032 583390 3088
rect 583446 3032 583451 3088
rect 350460 3030 583451 3032
rect 350460 3028 350466 3030
rect 583385 3027 583451 3030
rect 223614 2954 223620 2956
rect 110505 2952 117882 2954
rect 110505 2896 110510 2952
rect 110566 2896 117882 2952
rect 110505 2894 117882 2896
rect 118006 2894 223620 2954
rect 106917 2891 106983 2894
rect 110505 2891 110571 2894
rect 60825 2818 60891 2821
rect 62062 2818 62068 2820
rect 60825 2816 62068 2818
rect 60825 2760 60830 2816
rect 60886 2760 62068 2816
rect 60825 2758 62068 2760
rect 60825 2755 60891 2758
rect 62062 2756 62068 2758
rect 62132 2756 62138 2820
rect 66713 2818 66779 2821
rect 71589 2818 71655 2821
rect 66713 2816 71655 2818
rect 66713 2760 66718 2816
rect 66774 2760 71594 2816
rect 71650 2760 71655 2816
rect 66713 2758 71655 2760
rect 66713 2755 66779 2758
rect 71589 2755 71655 2758
rect 92749 2818 92815 2821
rect 115974 2818 115980 2820
rect 92749 2816 115980 2818
rect 92749 2760 92754 2816
rect 92810 2760 115980 2816
rect 92749 2758 115980 2760
rect 92749 2755 92815 2758
rect 115974 2756 115980 2758
rect 116044 2756 116050 2820
rect 117822 2818 117882 2894
rect 223614 2892 223620 2894
rect 223684 2892 223690 2956
rect 360193 2954 360259 2957
rect 360694 2954 360700 2956
rect 360193 2952 360700 2954
rect 360193 2896 360198 2952
rect 360254 2896 360700 2952
rect 360193 2894 360700 2896
rect 360193 2891 360259 2894
rect 360694 2892 360700 2894
rect 360764 2892 360770 2956
rect 376753 2954 376819 2957
rect 377254 2954 377260 2956
rect 376753 2952 377260 2954
rect 376753 2896 376758 2952
rect 376814 2896 377260 2952
rect 376753 2894 377260 2896
rect 376753 2891 376819 2894
rect 377254 2892 377260 2894
rect 377324 2892 377330 2956
rect 127014 2818 127020 2820
rect 117822 2758 127020 2818
rect 127014 2756 127020 2758
rect 127084 2756 127090 2820
<< via3 >>
rect 219204 699756 219268 699820
rect 251772 543628 251836 543692
rect 277900 543492 277964 543556
rect 327580 543356 327644 543420
rect 228220 543220 228284 543284
rect 230980 543084 231044 543148
rect 255820 543084 255884 543148
rect 280660 542948 280724 543012
rect 331812 542948 331876 543012
rect 335860 542948 335924 543012
rect 271092 542812 271156 542876
rect 322060 542812 322124 542876
rect 363460 542812 363524 542876
rect 197860 542676 197924 542740
rect 367692 542676 367756 542740
rect 137140 542540 137204 542604
rect 166212 542540 166276 542604
rect 222700 542540 222764 542604
rect 242020 542540 242084 542604
rect 266860 542540 266924 542604
rect 353892 542540 353956 542604
rect 389772 542540 389836 542604
rect 152412 542404 152476 542468
rect 161980 542404 162044 542468
rect 208900 542404 208964 542468
rect 237972 542404 238036 542468
rect 250300 542404 250364 542468
rect 304948 541044 305012 541108
rect 72924 539548 72988 539612
rect 75684 539608 75748 539612
rect 75684 539552 75698 539608
rect 75698 539552 75748 539608
rect 75684 539548 75748 539552
rect 106780 539548 106844 539612
rect 115980 539548 116044 539612
rect 119844 539548 119908 539612
rect 125364 539608 125428 539612
rect 125364 539552 125378 539608
rect 125378 539552 125428 539608
rect 125364 539548 125428 539552
rect 127020 539548 127084 539612
rect 155724 539548 155788 539612
rect 219940 539548 220004 539612
rect 246252 539548 246316 539612
rect 252508 539548 252572 539612
rect 283788 539608 283852 539612
rect 283788 539552 283838 539608
rect 283838 539552 283852 539608
rect 283788 539548 283852 539552
rect 313228 539548 313292 539612
rect 330340 539548 330404 539612
rect 341196 539548 341260 539612
rect 360700 539548 360764 539612
rect 377260 539608 377324 539612
rect 377260 539552 377310 539608
rect 377310 539552 377324 539608
rect 377260 539548 377324 539552
rect 382228 539548 382292 539612
rect 384988 539548 385052 539612
rect 387932 539548 387996 539612
rect 393820 539548 393884 539612
rect 400812 539548 400876 539612
rect 223620 539412 223684 539476
rect 240364 539412 240428 539476
rect 269620 539412 269684 539476
rect 279004 539412 279068 539476
rect 298140 539472 298204 539476
rect 298140 539416 298190 539472
rect 298190 539416 298204 539472
rect 298140 539412 298204 539416
rect 309180 539472 309244 539476
rect 309180 539416 309194 539472
rect 309194 539416 309244 539472
rect 309180 539412 309244 539416
rect 350396 539472 350460 539476
rect 350396 539416 350410 539472
rect 350410 539416 350460 539472
rect 350396 539412 350460 539416
rect 439452 488548 439516 488612
rect 60596 485828 60660 485892
rect 33732 462300 33796 462364
rect 439452 433468 439516 433532
rect 439268 425716 439332 425780
rect 453252 418236 453316 418300
rect 450492 404364 450556 404428
rect 21220 398652 21284 398716
rect 439452 398108 439516 398172
rect 439452 392668 439516 392732
rect 500172 378116 500236 378180
rect 60596 370636 60660 370700
rect 439452 347244 439516 347308
rect 60596 343708 60660 343772
rect 471100 311884 471164 311948
rect 35020 306308 35084 306372
rect 60596 303316 60660 303380
rect 439452 302092 439516 302156
rect 449940 302092 450004 302156
rect 449940 298148 450004 298212
rect 60596 274484 60660 274548
rect 450492 231916 450556 231980
rect 60596 213148 60660 213212
rect 36492 202812 36556 202876
rect 60596 179284 60660 179348
rect 60596 160788 60660 160852
rect 453252 138076 453316 138140
rect 468340 125564 468404 125628
rect 32260 111692 32324 111756
rect 22692 97820 22756 97884
rect 219204 57836 219268 57900
rect 367692 40564 367756 40628
rect 152412 26828 152476 26892
rect 219940 24108 220004 24172
rect 388116 24108 388180 24172
rect 269620 21388 269684 21452
rect 161980 21252 162044 21316
rect 251772 21252 251836 21316
rect 384988 18668 385052 18732
rect 119844 18532 119908 18596
rect 240364 17444 240428 17508
rect 155724 17308 155788 17372
rect 125364 17172 125428 17236
rect 222700 15812 222764 15876
rect 313228 15812 313292 15876
rect 353892 15812 353956 15876
rect 363460 14588 363524 14652
rect 106780 14452 106844 14516
rect 208900 13092 208964 13156
rect 400812 12956 400876 13020
rect 242020 12004 242084 12068
rect 166212 11868 166276 11932
rect 228220 11732 228284 11796
rect 237972 11732 238036 11796
rect 322060 11596 322124 11660
rect 255820 10916 255884 10980
rect 280660 10372 280724 10436
rect 327580 10372 327644 10436
rect 246252 10236 246316 10300
rect 341196 9556 341260 9620
rect 389772 9012 389836 9076
rect 382228 8876 382292 8940
rect 137140 7652 137204 7716
rect 250300 5612 250364 5676
rect 266860 5612 266924 5676
rect 335860 5612 335924 5676
rect 197860 4116 197924 4180
rect 230980 4116 231044 4180
rect 271092 4116 271156 4180
rect 277900 4116 277964 4180
rect 331812 4116 331876 4180
rect 72924 3980 72988 4044
rect 298140 3980 298204 4044
rect 393820 3980 393884 4044
rect 252508 3164 252572 3228
rect 279004 3164 279068 3228
rect 75684 3028 75748 3092
rect 283788 3028 283852 3092
rect 304948 3028 305012 3092
rect 330340 3028 330404 3092
rect 350396 3028 350460 3092
rect 62068 2756 62132 2820
rect 115980 2756 116044 2820
rect 223620 2892 223684 2956
rect 360700 2892 360764 2956
rect 377260 2892 377324 2956
rect 127020 2756 127084 2820
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 21222 398717 21282 425902
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 21219 398716 21285 398717
rect 21219 398652 21220 398716
rect 21284 398652 21285 398716
rect 21219 398651 21285 398652
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 22694 97885 22754 397342
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 22691 97884 22757 97885
rect 22691 97820 22692 97884
rect 22756 97820 22757 97884
rect 22691 97819 22757 97820
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 33731 462364 33797 462365
rect 33731 462300 33732 462364
rect 33796 462300 33797 462364
rect 33731 462299 33797 462300
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 32262 111757 32322 391222
rect 33734 347258 33794 462299
rect 35022 306373 35082 487782
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 35019 306372 35085 306373
rect 35019 306308 35020 306372
rect 35084 306308 35085 306372
rect 35019 306307 35085 306308
rect 36494 202877 36554 433382
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 36491 202876 36557 202877
rect 36491 202812 36492 202876
rect 36556 202812 36557 202876
rect 36491 202811 36557 202812
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 32259 111756 32325 111757
rect 32259 111692 32260 111756
rect 32324 111692 32325 111756
rect 32259 111691 32325 111692
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 542000 60134 564618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 542000 63854 568338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 542000 67574 572058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 542000 74414 542898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 542000 78134 546618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 542000 81854 550338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 542000 85574 554058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 542000 92414 560898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 542000 96134 564618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 542000 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 542000 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 542000 110414 542898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 542000 114134 546618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 542000 117854 550338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 542000 121574 554058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 542000 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 542000 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 542000 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 137139 542604 137205 542605
rect 137139 542540 137140 542604
rect 137204 542540 137205 542604
rect 137139 542539 137205 542540
rect 72923 539612 72989 539613
rect 72923 539548 72924 539612
rect 72988 539548 72989 539612
rect 72923 539547 72989 539548
rect 75683 539612 75749 539613
rect 75683 539548 75684 539612
rect 75748 539548 75749 539612
rect 75683 539547 75749 539548
rect 106779 539612 106845 539613
rect 106779 539548 106780 539612
rect 106844 539548 106845 539612
rect 106779 539547 106845 539548
rect 115979 539612 116045 539613
rect 115979 539548 115980 539612
rect 116044 539548 116045 539612
rect 115979 539547 116045 539548
rect 119843 539612 119909 539613
rect 119843 539548 119844 539612
rect 119908 539548 119909 539612
rect 119843 539547 119909 539548
rect 125363 539612 125429 539613
rect 125363 539548 125364 539612
rect 125428 539548 125429 539612
rect 125363 539547 125429 539548
rect 127019 539612 127085 539613
rect 127019 539548 127020 539612
rect 127084 539548 127085 539612
rect 127019 539547 127085 539548
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 64208 471454 64528 471486
rect 64208 471218 64250 471454
rect 64486 471218 64528 471454
rect 64208 471134 64528 471218
rect 64208 470898 64250 471134
rect 64486 470898 64528 471134
rect 64208 470866 64528 470898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 64208 435454 64528 435486
rect 64208 435218 64250 435454
rect 64486 435218 64528 435454
rect 64208 435134 64528 435218
rect 64208 434898 64250 435134
rect 64486 434898 64528 435134
rect 64208 434866 64528 434898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 64208 399454 64528 399486
rect 64208 399218 64250 399454
rect 64486 399218 64528 399454
rect 64208 399134 64528 399218
rect 64208 398898 64250 399134
rect 64486 398898 64528 399134
rect 64208 398866 64528 398898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 60598 370701 60658 371502
rect 60595 370700 60661 370701
rect 60595 370636 60596 370700
rect 60660 370636 60661 370700
rect 60595 370635 60661 370636
rect 64208 363454 64528 363486
rect 64208 363218 64250 363454
rect 64486 363218 64528 363454
rect 64208 363134 64528 363218
rect 64208 362898 64250 363134
rect 64486 362898 64528 363134
rect 64208 362866 64528 362898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 64208 327454 64528 327486
rect 64208 327218 64250 327454
rect 64486 327218 64528 327454
rect 64208 327134 64528 327218
rect 64208 326898 64250 327134
rect 64486 326898 64528 327134
rect 64208 326866 64528 326898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 60598 303381 60658 303502
rect 60595 303380 60661 303381
rect 60595 303316 60596 303380
rect 60660 303316 60661 303380
rect 60595 303315 60661 303316
rect 65382 301018 65442 303502
rect 64208 291454 64528 291486
rect 64208 291218 64250 291454
rect 64486 291218 64528 291454
rect 64208 291134 64528 291218
rect 64208 290898 64250 291134
rect 64486 290898 64528 291134
rect 64208 290866 64528 290898
rect 60595 274548 60661 274549
rect 60595 274498 60596 274548
rect 60660 274498 60661 274548
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 64208 255454 64528 255486
rect 64208 255218 64250 255454
rect 64486 255218 64528 255454
rect 64208 255134 64528 255218
rect 64208 254898 64250 255134
rect 64486 254898 64528 255134
rect 64208 254866 64528 254898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 64208 219454 64528 219486
rect 64208 219218 64250 219454
rect 64486 219218 64528 219454
rect 64208 219134 64528 219218
rect 64208 218898 64250 219134
rect 64486 218898 64528 219134
rect 64208 218866 64528 218898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 64208 183454 64528 183486
rect 64208 183218 64250 183454
rect 64486 183218 64528 183454
rect 64208 183134 64528 183218
rect 64208 182898 64250 183134
rect 64486 182898 64528 183134
rect 64208 182866 64528 182898
rect 60595 179348 60661 179349
rect 60595 179298 60596 179348
rect 60660 179298 60661 179348
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 64208 111454 64528 111486
rect 64208 111218 64250 111454
rect 64486 111218 64528 111454
rect 64208 111134 64528 111218
rect 64208 110898 64250 111134
rect 64486 110898 64528 111134
rect 64208 110866 64528 110898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 64208 75454 64528 75486
rect 64208 75218 64250 75454
rect 64486 75218 64528 75454
rect 64208 75134 64528 75218
rect 64208 74898 64250 75134
rect 64486 74898 64528 75134
rect 64208 74866 64528 74898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 62070 2821 62130 4302
rect 62067 2820 62133 2821
rect 62067 2756 62068 2820
rect 62132 2756 62133 2820
rect 62067 2755 62133 2756
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 72926 4045 72986 539547
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 72923 4044 72989 4045
rect 72923 3980 72924 4044
rect 72988 3980 72989 4044
rect 72923 3979 72989 3980
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 75686 3093 75746 539547
rect 79568 525454 79888 525486
rect 79568 525218 79610 525454
rect 79846 525218 79888 525454
rect 79568 525134 79888 525218
rect 79568 524898 79610 525134
rect 79846 524898 79888 525134
rect 79568 524866 79888 524898
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 79568 489454 79888 489486
rect 79568 489218 79610 489454
rect 79846 489218 79888 489454
rect 79568 489134 79888 489218
rect 79568 488898 79610 489134
rect 79846 488898 79888 489134
rect 79568 488866 79888 488898
rect 94928 471454 95248 471486
rect 94928 471218 94970 471454
rect 95206 471218 95248 471454
rect 94928 471134 95248 471218
rect 94928 470898 94970 471134
rect 95206 470898 95248 471134
rect 94928 470866 95248 470898
rect 79568 453454 79888 453486
rect 79568 453218 79610 453454
rect 79846 453218 79888 453454
rect 79568 453134 79888 453218
rect 79568 452898 79610 453134
rect 79846 452898 79888 453134
rect 79568 452866 79888 452898
rect 94928 435454 95248 435486
rect 94928 435218 94970 435454
rect 95206 435218 95248 435454
rect 94928 435134 95248 435218
rect 94928 434898 94970 435134
rect 95206 434898 95248 435134
rect 94928 434866 95248 434898
rect 79568 417454 79888 417486
rect 79568 417218 79610 417454
rect 79846 417218 79888 417454
rect 79568 417134 79888 417218
rect 79568 416898 79610 417134
rect 79846 416898 79888 417134
rect 79568 416866 79888 416898
rect 94928 399454 95248 399486
rect 94928 399218 94970 399454
rect 95206 399218 95248 399454
rect 94928 399134 95248 399218
rect 94928 398898 94970 399134
rect 95206 398898 95248 399134
rect 94928 398866 95248 398898
rect 79568 381454 79888 381486
rect 79568 381218 79610 381454
rect 79846 381218 79888 381454
rect 79568 381134 79888 381218
rect 79568 380898 79610 381134
rect 79846 380898 79888 381134
rect 79568 380866 79888 380898
rect 94928 363454 95248 363486
rect 94928 363218 94970 363454
rect 95206 363218 95248 363454
rect 94928 363134 95248 363218
rect 94928 362898 94970 363134
rect 95206 362898 95248 363134
rect 94928 362866 95248 362898
rect 79568 345454 79888 345486
rect 79568 345218 79610 345454
rect 79846 345218 79888 345454
rect 79568 345134 79888 345218
rect 79568 344898 79610 345134
rect 79846 344898 79888 345134
rect 79568 344866 79888 344898
rect 94928 327454 95248 327486
rect 94928 327218 94970 327454
rect 95206 327218 95248 327454
rect 94928 327134 95248 327218
rect 94928 326898 94970 327134
rect 95206 326898 95248 327134
rect 94928 326866 95248 326898
rect 79568 309454 79888 309486
rect 79568 309218 79610 309454
rect 79846 309218 79888 309454
rect 79568 309134 79888 309218
rect 79568 308898 79610 309134
rect 79846 308898 79888 309134
rect 79568 308866 79888 308898
rect 85438 301018 85498 303502
rect 93902 301018 93962 303502
rect 94928 291454 95248 291486
rect 94928 291218 94970 291454
rect 95206 291218 95248 291454
rect 94928 291134 95248 291218
rect 94928 290898 94970 291134
rect 95206 290898 95248 291134
rect 94928 290866 95248 290898
rect 79568 273454 79888 273486
rect 79568 273218 79610 273454
rect 79846 273218 79888 273454
rect 79568 273134 79888 273218
rect 79568 272898 79610 273134
rect 79846 272898 79888 273134
rect 79568 272866 79888 272898
rect 94928 255454 95248 255486
rect 94928 255218 94970 255454
rect 95206 255218 95248 255454
rect 94928 255134 95248 255218
rect 94928 254898 94970 255134
rect 95206 254898 95248 255134
rect 94928 254866 95248 254898
rect 79568 237454 79888 237486
rect 79568 237218 79610 237454
rect 79846 237218 79888 237454
rect 79568 237134 79888 237218
rect 79568 236898 79610 237134
rect 79846 236898 79888 237134
rect 79568 236866 79888 236898
rect 94928 219454 95248 219486
rect 94928 219218 94970 219454
rect 95206 219218 95248 219454
rect 94928 219134 95248 219218
rect 94928 218898 94970 219134
rect 95206 218898 95248 219134
rect 94928 218866 95248 218898
rect 79568 201454 79888 201486
rect 79568 201218 79610 201454
rect 79846 201218 79888 201454
rect 79568 201134 79888 201218
rect 79568 200898 79610 201134
rect 79846 200898 79888 201134
rect 79568 200866 79888 200898
rect 94928 183454 95248 183486
rect 94928 183218 94970 183454
rect 95206 183218 95248 183454
rect 94928 183134 95248 183218
rect 94928 182898 94970 183134
rect 95206 182898 95248 183134
rect 94928 182866 95248 182898
rect 79568 165454 79888 165486
rect 79568 165218 79610 165454
rect 79846 165218 79888 165454
rect 79568 165134 79888 165218
rect 79568 164898 79610 165134
rect 79846 164898 79888 165134
rect 79568 164866 79888 164898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 79568 129454 79888 129486
rect 79568 129218 79610 129454
rect 79846 129218 79888 129454
rect 79568 129134 79888 129218
rect 79568 128898 79610 129134
rect 79846 128898 79888 129134
rect 79568 128866 79888 128898
rect 94928 111454 95248 111486
rect 94928 111218 94970 111454
rect 95206 111218 95248 111454
rect 94928 111134 95248 111218
rect 94928 110898 94970 111134
rect 95206 110898 95248 111134
rect 94928 110866 95248 110898
rect 79568 93454 79888 93486
rect 79568 93218 79610 93454
rect 79846 93218 79888 93454
rect 79568 93134 79888 93218
rect 79568 92898 79610 93134
rect 79846 92898 79888 93134
rect 79568 92866 79888 92898
rect 94928 75454 95248 75486
rect 94928 75218 94970 75454
rect 95206 75218 95248 75454
rect 94928 75134 95248 75218
rect 94928 74898 94970 75134
rect 95206 74898 95248 75134
rect 94928 74866 95248 74898
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 75683 3092 75749 3093
rect 75683 3028 75684 3092
rect 75748 3028 75749 3092
rect 75683 3027 75749 3028
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 106782 14517 106842 539547
rect 110288 525454 110608 525486
rect 110288 525218 110330 525454
rect 110566 525218 110608 525454
rect 110288 525134 110608 525218
rect 110288 524898 110330 525134
rect 110566 524898 110608 525134
rect 110288 524866 110608 524898
rect 110288 489454 110608 489486
rect 110288 489218 110330 489454
rect 110566 489218 110608 489454
rect 110288 489134 110608 489218
rect 110288 488898 110330 489134
rect 110566 488898 110608 489134
rect 110288 488866 110608 488898
rect 110288 453454 110608 453486
rect 110288 453218 110330 453454
rect 110566 453218 110608 453454
rect 110288 453134 110608 453218
rect 110288 452898 110330 453134
rect 110566 452898 110608 453134
rect 110288 452866 110608 452898
rect 110288 417454 110608 417486
rect 110288 417218 110330 417454
rect 110566 417218 110608 417454
rect 110288 417134 110608 417218
rect 110288 416898 110330 417134
rect 110566 416898 110608 417134
rect 110288 416866 110608 416898
rect 110288 381454 110608 381486
rect 110288 381218 110330 381454
rect 110566 381218 110608 381454
rect 110288 381134 110608 381218
rect 110288 380898 110330 381134
rect 110566 380898 110608 381134
rect 110288 380866 110608 380898
rect 110288 345454 110608 345486
rect 110288 345218 110330 345454
rect 110566 345218 110608 345454
rect 110288 345134 110608 345218
rect 110288 344898 110330 345134
rect 110566 344898 110608 345134
rect 110288 344866 110608 344898
rect 115982 325710 116042 539547
rect 115982 325650 116410 325710
rect 110288 309454 110608 309486
rect 110288 309218 110330 309454
rect 110566 309218 110608 309454
rect 110288 309134 110608 309218
rect 110288 308898 110330 309134
rect 110566 308898 110608 309134
rect 110288 308866 110608 308898
rect 113774 301018 113834 303502
rect 116350 296730 116410 325650
rect 115982 296670 116410 296730
rect 110288 273454 110608 273486
rect 110288 273218 110330 273454
rect 110566 273218 110608 273454
rect 110288 273134 110608 273218
rect 110288 272898 110330 273134
rect 110566 272898 110608 273134
rect 110288 272866 110608 272898
rect 110288 237454 110608 237486
rect 110288 237218 110330 237454
rect 110566 237218 110608 237454
rect 110288 237134 110608 237218
rect 110288 236898 110330 237134
rect 110566 236898 110608 237134
rect 110288 236866 110608 236898
rect 110288 201454 110608 201486
rect 110288 201218 110330 201454
rect 110566 201218 110608 201454
rect 110288 201134 110608 201218
rect 110288 200898 110330 201134
rect 110566 200898 110608 201134
rect 110288 200866 110608 200898
rect 110288 165454 110608 165486
rect 110288 165218 110330 165454
rect 110566 165218 110608 165454
rect 110288 165134 110608 165218
rect 110288 164898 110330 165134
rect 110566 164898 110608 165134
rect 110288 164866 110608 164898
rect 110288 129454 110608 129486
rect 110288 129218 110330 129454
rect 110566 129218 110608 129454
rect 110288 129134 110608 129218
rect 110288 128898 110330 129134
rect 110566 128898 110608 129134
rect 110288 128866 110608 128898
rect 110288 93454 110608 93486
rect 110288 93218 110330 93454
rect 110566 93218 110608 93454
rect 110288 93134 110608 93218
rect 110288 92898 110330 93134
rect 110566 92898 110608 93134
rect 110288 92866 110608 92898
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 106779 14516 106845 14517
rect 106779 14452 106780 14516
rect 106844 14452 106845 14516
rect 106779 14451 106845 14452
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 115982 2821 116042 296670
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 119846 18597 119906 539547
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 119843 18596 119909 18597
rect 119843 18532 119844 18596
rect 119908 18532 119909 18596
rect 119843 18531 119909 18532
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 115979 2820 116045 2821
rect 115979 2756 115980 2820
rect 116044 2756 116045 2820
rect 115979 2755 116045 2756
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 14614 121574 50058
rect 125366 17237 125426 539547
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 125648 471454 125968 471486
rect 125648 471218 125690 471454
rect 125926 471218 125968 471454
rect 125648 471134 125968 471218
rect 125648 470898 125690 471134
rect 125926 470898 125968 471134
rect 125648 470866 125968 470898
rect 125648 435454 125968 435486
rect 125648 435218 125690 435454
rect 125926 435218 125968 435454
rect 125648 435134 125968 435218
rect 125648 434898 125690 435134
rect 125926 434898 125968 435134
rect 125648 434866 125968 434898
rect 125648 399454 125968 399486
rect 125648 399218 125690 399454
rect 125926 399218 125968 399454
rect 125648 399134 125968 399218
rect 125648 398898 125690 399134
rect 125926 398898 125968 399134
rect 125648 398866 125968 398898
rect 125648 363454 125968 363486
rect 125648 363218 125690 363454
rect 125926 363218 125968 363454
rect 125648 363134 125968 363218
rect 125648 362898 125690 363134
rect 125926 362898 125968 363134
rect 125648 362866 125968 362898
rect 125648 327454 125968 327486
rect 125648 327218 125690 327454
rect 125926 327218 125968 327454
rect 125648 327134 125968 327218
rect 125648 326898 125690 327134
rect 125926 326898 125968 327134
rect 125648 326866 125968 326898
rect 125648 291454 125968 291486
rect 125648 291218 125690 291454
rect 125926 291218 125968 291454
rect 125648 291134 125968 291218
rect 125648 290898 125690 291134
rect 125926 290898 125968 291134
rect 125648 290866 125968 290898
rect 125648 255454 125968 255486
rect 125648 255218 125690 255454
rect 125926 255218 125968 255454
rect 125648 255134 125968 255218
rect 125648 254898 125690 255134
rect 125926 254898 125968 255134
rect 125648 254866 125968 254898
rect 125648 219454 125968 219486
rect 125648 219218 125690 219454
rect 125926 219218 125968 219454
rect 125648 219134 125968 219218
rect 125648 218898 125690 219134
rect 125926 218898 125968 219134
rect 125648 218866 125968 218898
rect 125648 183454 125968 183486
rect 125648 183218 125690 183454
rect 125926 183218 125968 183454
rect 125648 183134 125968 183218
rect 125648 182898 125690 183134
rect 125926 182898 125968 183134
rect 125648 182866 125968 182898
rect 125648 147454 125968 147486
rect 125648 147218 125690 147454
rect 125926 147218 125968 147454
rect 125648 147134 125968 147218
rect 125648 146898 125690 147134
rect 125926 146898 125968 147134
rect 125648 146866 125968 146898
rect 125648 111454 125968 111486
rect 125648 111218 125690 111454
rect 125926 111218 125968 111454
rect 125648 111134 125968 111218
rect 125648 110898 125690 111134
rect 125926 110898 125968 111134
rect 125648 110866 125968 110898
rect 125648 75454 125968 75486
rect 125648 75218 125690 75454
rect 125926 75218 125968 75454
rect 125648 75134 125968 75218
rect 125648 74898 125690 75134
rect 125926 74898 125968 75134
rect 125648 74866 125968 74898
rect 125363 17236 125429 17237
rect 125363 17172 125364 17236
rect 125428 17172 125429 17236
rect 125363 17171 125429 17172
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127022 2821 127082 539547
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127019 2820 127085 2821
rect 127019 2756 127020 2820
rect 127084 2756 127085 2820
rect 127019 2755 127085 2756
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 137142 7717 137202 542539
rect 138954 542000 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 542000 146414 542898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 542000 150134 546618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 152411 542468 152477 542469
rect 152411 542404 152412 542468
rect 152476 542404 152477 542468
rect 152411 542403 152477 542404
rect 141008 525454 141328 525486
rect 141008 525218 141050 525454
rect 141286 525218 141328 525454
rect 141008 525134 141328 525218
rect 141008 524898 141050 525134
rect 141286 524898 141328 525134
rect 141008 524866 141328 524898
rect 141008 489454 141328 489486
rect 141008 489218 141050 489454
rect 141286 489218 141328 489454
rect 141008 489134 141328 489218
rect 141008 488898 141050 489134
rect 141286 488898 141328 489134
rect 141008 488866 141328 488898
rect 141008 453454 141328 453486
rect 141008 453218 141050 453454
rect 141286 453218 141328 453454
rect 141008 453134 141328 453218
rect 141008 452898 141050 453134
rect 141286 452898 141328 453134
rect 141008 452866 141328 452898
rect 141008 417454 141328 417486
rect 141008 417218 141050 417454
rect 141286 417218 141328 417454
rect 141008 417134 141328 417218
rect 141008 416898 141050 417134
rect 141286 416898 141328 417134
rect 141008 416866 141328 416898
rect 141008 381454 141328 381486
rect 141008 381218 141050 381454
rect 141286 381218 141328 381454
rect 141008 381134 141328 381218
rect 141008 380898 141050 381134
rect 141286 380898 141328 381134
rect 141008 380866 141328 380898
rect 141008 345454 141328 345486
rect 141008 345218 141050 345454
rect 141286 345218 141328 345454
rect 141008 345134 141328 345218
rect 141008 344898 141050 345134
rect 141286 344898 141328 345134
rect 141008 344866 141328 344898
rect 141008 309454 141328 309486
rect 141008 309218 141050 309454
rect 141286 309218 141328 309454
rect 141008 309134 141328 309218
rect 141008 308898 141050 309134
rect 141286 308898 141328 309134
rect 141008 308866 141328 308898
rect 143030 301018 143090 303502
rect 141008 273454 141328 273486
rect 141008 273218 141050 273454
rect 141286 273218 141328 273454
rect 141008 273134 141328 273218
rect 141008 272898 141050 273134
rect 141286 272898 141328 273134
rect 141008 272866 141328 272898
rect 141008 237454 141328 237486
rect 141008 237218 141050 237454
rect 141286 237218 141328 237454
rect 141008 237134 141328 237218
rect 141008 236898 141050 237134
rect 141286 236898 141328 237134
rect 141008 236866 141328 236898
rect 141008 201454 141328 201486
rect 141008 201218 141050 201454
rect 141286 201218 141328 201454
rect 141008 201134 141328 201218
rect 141008 200898 141050 201134
rect 141286 200898 141328 201134
rect 141008 200866 141328 200898
rect 141008 165454 141328 165486
rect 141008 165218 141050 165454
rect 141286 165218 141328 165454
rect 141008 165134 141328 165218
rect 141008 164898 141050 165134
rect 141286 164898 141328 165134
rect 141008 164866 141328 164898
rect 141008 129454 141328 129486
rect 141008 129218 141050 129454
rect 141286 129218 141328 129454
rect 141008 129134 141328 129218
rect 141008 128898 141050 129134
rect 141286 128898 141328 129134
rect 141008 128866 141328 128898
rect 141008 93454 141328 93486
rect 141008 93218 141050 93454
rect 141286 93218 141328 93454
rect 141008 93134 141328 93218
rect 141008 92898 141050 93134
rect 141286 92898 141328 93134
rect 141008 92866 141328 92898
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 137139 7716 137205 7717
rect 137139 7652 137140 7716
rect 137204 7652 137205 7716
rect 137139 7651 137205 7652
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 152414 26893 152474 542403
rect 153234 542000 153854 550338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 542000 157574 554058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 161979 542468 162045 542469
rect 161979 542404 161980 542468
rect 162044 542404 162045 542468
rect 161979 542403 162045 542404
rect 155723 539612 155789 539613
rect 155723 539548 155724 539612
rect 155788 539548 155789 539612
rect 155723 539547 155789 539548
rect 153886 301018 153946 303502
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 152411 26892 152477 26893
rect 152411 26828 152412 26892
rect 152476 26828 152477 26892
rect 152411 26827 152477 26828
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 46338
rect 155726 17373 155786 539547
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 156368 471454 156688 471486
rect 156368 471218 156410 471454
rect 156646 471218 156688 471454
rect 156368 471134 156688 471218
rect 156368 470898 156410 471134
rect 156646 470898 156688 471134
rect 156368 470866 156688 470898
rect 156368 435454 156688 435486
rect 156368 435218 156410 435454
rect 156646 435218 156688 435454
rect 156368 435134 156688 435218
rect 156368 434898 156410 435134
rect 156646 434898 156688 435134
rect 156368 434866 156688 434898
rect 156368 399454 156688 399486
rect 156368 399218 156410 399454
rect 156646 399218 156688 399454
rect 156368 399134 156688 399218
rect 156368 398898 156410 399134
rect 156646 398898 156688 399134
rect 156368 398866 156688 398898
rect 156368 363454 156688 363486
rect 156368 363218 156410 363454
rect 156646 363218 156688 363454
rect 156368 363134 156688 363218
rect 156368 362898 156410 363134
rect 156646 362898 156688 363134
rect 156368 362866 156688 362898
rect 156368 327454 156688 327486
rect 156368 327218 156410 327454
rect 156646 327218 156688 327454
rect 156368 327134 156688 327218
rect 156368 326898 156410 327134
rect 156646 326898 156688 327134
rect 156368 326866 156688 326898
rect 161614 301018 161674 303502
rect 156368 291454 156688 291486
rect 156368 291218 156410 291454
rect 156646 291218 156688 291454
rect 156368 291134 156688 291218
rect 156368 290898 156410 291134
rect 156646 290898 156688 291134
rect 156368 290866 156688 290898
rect 156368 255454 156688 255486
rect 156368 255218 156410 255454
rect 156646 255218 156688 255454
rect 156368 255134 156688 255218
rect 156368 254898 156410 255134
rect 156646 254898 156688 255134
rect 156368 254866 156688 254898
rect 156368 219454 156688 219486
rect 156368 219218 156410 219454
rect 156646 219218 156688 219454
rect 156368 219134 156688 219218
rect 156368 218898 156410 219134
rect 156646 218898 156688 219134
rect 156368 218866 156688 218898
rect 156368 183454 156688 183486
rect 156368 183218 156410 183454
rect 156646 183218 156688 183454
rect 156368 183134 156688 183218
rect 156368 182898 156410 183134
rect 156646 182898 156688 183134
rect 156368 182866 156688 182898
rect 156368 147454 156688 147486
rect 156368 147218 156410 147454
rect 156646 147218 156688 147454
rect 156368 147134 156688 147218
rect 156368 146898 156410 147134
rect 156646 146898 156688 147134
rect 156368 146866 156688 146898
rect 156368 111454 156688 111486
rect 156368 111218 156410 111454
rect 156646 111218 156688 111454
rect 156368 111134 156688 111218
rect 156368 110898 156410 111134
rect 156646 110898 156688 111134
rect 156368 110866 156688 110898
rect 156368 75454 156688 75486
rect 156368 75218 156410 75454
rect 156646 75218 156688 75454
rect 156368 75134 156688 75218
rect 156368 74898 156410 75134
rect 156646 74898 156688 75134
rect 156368 74866 156688 74898
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 155723 17372 155789 17373
rect 155723 17308 155724 17372
rect 155788 17308 155789 17372
rect 155723 17307 155789 17308
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 14614 157574 50058
rect 161982 21317 162042 542403
rect 163794 542000 164414 560898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 166211 542604 166277 542605
rect 166211 542540 166212 542604
rect 166276 542540 166277 542604
rect 166211 542539 166277 542540
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 161979 21316 162045 21317
rect 161979 21252 161980 21316
rect 162044 21252 162045 21316
rect 161979 21251 162045 21252
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 166214 11933 166274 542539
rect 167514 542000 168134 564618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 542000 171854 568338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 542000 175574 572058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 542000 182414 542898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 542000 186134 546618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 542000 189854 550338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 542000 193574 554058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 197859 542740 197925 542741
rect 197859 542676 197860 542740
rect 197924 542676 197925 542740
rect 197859 542675 197925 542676
rect 171728 525454 172048 525486
rect 171728 525218 171770 525454
rect 172006 525218 172048 525454
rect 171728 525134 172048 525218
rect 171728 524898 171770 525134
rect 172006 524898 172048 525134
rect 171728 524866 172048 524898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 171728 489454 172048 489486
rect 171728 489218 171770 489454
rect 172006 489218 172048 489454
rect 171728 489134 172048 489218
rect 171728 488898 171770 489134
rect 172006 488898 172048 489134
rect 171728 488866 172048 488898
rect 187088 471454 187408 471486
rect 187088 471218 187130 471454
rect 187366 471218 187408 471454
rect 187088 471134 187408 471218
rect 187088 470898 187130 471134
rect 187366 470898 187408 471134
rect 187088 470866 187408 470898
rect 171728 453454 172048 453486
rect 171728 453218 171770 453454
rect 172006 453218 172048 453454
rect 171728 453134 172048 453218
rect 171728 452898 171770 453134
rect 172006 452898 172048 453134
rect 171728 452866 172048 452898
rect 187088 435454 187408 435486
rect 187088 435218 187130 435454
rect 187366 435218 187408 435454
rect 187088 435134 187408 435218
rect 187088 434898 187130 435134
rect 187366 434898 187408 435134
rect 187088 434866 187408 434898
rect 171728 417454 172048 417486
rect 171728 417218 171770 417454
rect 172006 417218 172048 417454
rect 171728 417134 172048 417218
rect 171728 416898 171770 417134
rect 172006 416898 172048 417134
rect 171728 416866 172048 416898
rect 187088 399454 187408 399486
rect 187088 399218 187130 399454
rect 187366 399218 187408 399454
rect 187088 399134 187408 399218
rect 187088 398898 187130 399134
rect 187366 398898 187408 399134
rect 187088 398866 187408 398898
rect 171728 381454 172048 381486
rect 171728 381218 171770 381454
rect 172006 381218 172048 381454
rect 171728 381134 172048 381218
rect 171728 380898 171770 381134
rect 172006 380898 172048 381134
rect 171728 380866 172048 380898
rect 187088 363454 187408 363486
rect 187088 363218 187130 363454
rect 187366 363218 187408 363454
rect 187088 363134 187408 363218
rect 187088 362898 187130 363134
rect 187366 362898 187408 363134
rect 187088 362866 187408 362898
rect 171728 345454 172048 345486
rect 171728 345218 171770 345454
rect 172006 345218 172048 345454
rect 171728 345134 172048 345218
rect 171728 344898 171770 345134
rect 172006 344898 172048 345134
rect 171728 344866 172048 344898
rect 187088 327454 187408 327486
rect 187088 327218 187130 327454
rect 187366 327218 187408 327454
rect 187088 327134 187408 327218
rect 187088 326898 187130 327134
rect 187366 326898 187408 327134
rect 187088 326866 187408 326898
rect 171728 309454 172048 309486
rect 171728 309218 171770 309454
rect 172006 309218 172048 309454
rect 171728 309134 172048 309218
rect 171728 308898 171770 309134
rect 172006 308898 172048 309134
rect 171728 308866 172048 308898
rect 190686 301018 190746 303502
rect 187088 291454 187408 291486
rect 187088 291218 187130 291454
rect 187366 291218 187408 291454
rect 187088 291134 187408 291218
rect 187088 290898 187130 291134
rect 187366 290898 187408 291134
rect 187088 290866 187408 290898
rect 171728 273454 172048 273486
rect 171728 273218 171770 273454
rect 172006 273218 172048 273454
rect 171728 273134 172048 273218
rect 171728 272898 171770 273134
rect 172006 272898 172048 273134
rect 171728 272866 172048 272898
rect 187088 255454 187408 255486
rect 187088 255218 187130 255454
rect 187366 255218 187408 255454
rect 187088 255134 187408 255218
rect 187088 254898 187130 255134
rect 187366 254898 187408 255134
rect 187088 254866 187408 254898
rect 171728 237454 172048 237486
rect 171728 237218 171770 237454
rect 172006 237218 172048 237454
rect 171728 237134 172048 237218
rect 171728 236898 171770 237134
rect 172006 236898 172048 237134
rect 171728 236866 172048 236898
rect 187088 219454 187408 219486
rect 187088 219218 187130 219454
rect 187366 219218 187408 219454
rect 187088 219134 187408 219218
rect 187088 218898 187130 219134
rect 187366 218898 187408 219134
rect 187088 218866 187408 218898
rect 171728 201454 172048 201486
rect 171728 201218 171770 201454
rect 172006 201218 172048 201454
rect 171728 201134 172048 201218
rect 171728 200898 171770 201134
rect 172006 200898 172048 201134
rect 171728 200866 172048 200898
rect 187088 183454 187408 183486
rect 187088 183218 187130 183454
rect 187366 183218 187408 183454
rect 187088 183134 187408 183218
rect 187088 182898 187130 183134
rect 187366 182898 187408 183134
rect 187088 182866 187408 182898
rect 171728 165454 172048 165486
rect 171728 165218 171770 165454
rect 172006 165218 172048 165454
rect 171728 165134 172048 165218
rect 171728 164898 171770 165134
rect 172006 164898 172048 165134
rect 171728 164866 172048 164898
rect 187088 147454 187408 147486
rect 187088 147218 187130 147454
rect 187366 147218 187408 147454
rect 187088 147134 187408 147218
rect 187088 146898 187130 147134
rect 187366 146898 187408 147134
rect 187088 146866 187408 146898
rect 171728 129454 172048 129486
rect 171728 129218 171770 129454
rect 172006 129218 172048 129454
rect 171728 129134 172048 129218
rect 171728 128898 171770 129134
rect 172006 128898 172048 129134
rect 171728 128866 172048 128898
rect 187088 111454 187408 111486
rect 187088 111218 187130 111454
rect 187366 111218 187408 111454
rect 187088 111134 187408 111218
rect 187088 110898 187130 111134
rect 187366 110898 187408 111134
rect 187088 110866 187408 110898
rect 171728 93454 172048 93486
rect 171728 93218 171770 93454
rect 172006 93218 172048 93454
rect 171728 93134 172048 93218
rect 171728 92898 171770 93134
rect 172006 92898 172048 93134
rect 171728 92866 172048 92898
rect 187088 75454 187408 75486
rect 187088 75218 187130 75454
rect 187366 75218 187408 75454
rect 187088 75134 187408 75218
rect 187088 74898 187130 75134
rect 187366 74898 187408 75134
rect 187088 74866 187408 74898
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 166211 11932 166277 11933
rect 166211 11868 166212 11932
rect 166276 11868 166277 11932
rect 166211 11867 166277 11868
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 197862 4181 197922 542675
rect 199794 542000 200414 560898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 542000 204134 564618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 542000 207854 568338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 208899 542468 208965 542469
rect 208899 542404 208900 542468
rect 208964 542404 208965 542468
rect 208899 542403 208965 542404
rect 202448 525454 202768 525486
rect 202448 525218 202490 525454
rect 202726 525218 202768 525454
rect 202448 525134 202768 525218
rect 202448 524898 202490 525134
rect 202726 524898 202768 525134
rect 202448 524866 202768 524898
rect 202448 489454 202768 489486
rect 202448 489218 202490 489454
rect 202726 489218 202768 489454
rect 202448 489134 202768 489218
rect 202448 488898 202490 489134
rect 202726 488898 202768 489134
rect 202448 488866 202768 488898
rect 202448 453454 202768 453486
rect 202448 453218 202490 453454
rect 202726 453218 202768 453454
rect 202448 453134 202768 453218
rect 202448 452898 202490 453134
rect 202726 452898 202768 453134
rect 202448 452866 202768 452898
rect 202448 417454 202768 417486
rect 202448 417218 202490 417454
rect 202726 417218 202768 417454
rect 202448 417134 202768 417218
rect 202448 416898 202490 417134
rect 202726 416898 202768 417134
rect 202448 416866 202768 416898
rect 202448 381454 202768 381486
rect 202448 381218 202490 381454
rect 202726 381218 202768 381454
rect 202448 381134 202768 381218
rect 202448 380898 202490 381134
rect 202726 380898 202768 381134
rect 202448 380866 202768 380898
rect 202448 345454 202768 345486
rect 202448 345218 202490 345454
rect 202726 345218 202768 345454
rect 202448 345134 202768 345218
rect 202448 344898 202490 345134
rect 202726 344898 202768 345134
rect 202448 344866 202768 344898
rect 202448 309454 202768 309486
rect 202448 309218 202490 309454
rect 202726 309218 202768 309454
rect 202448 309134 202768 309218
rect 202448 308898 202490 309134
rect 202726 308898 202768 309134
rect 202448 308866 202768 308898
rect 202448 273454 202768 273486
rect 202448 273218 202490 273454
rect 202726 273218 202768 273454
rect 202448 273134 202768 273218
rect 202448 272898 202490 273134
rect 202726 272898 202768 273134
rect 202448 272866 202768 272898
rect 202448 237454 202768 237486
rect 202448 237218 202490 237454
rect 202726 237218 202768 237454
rect 202448 237134 202768 237218
rect 202448 236898 202490 237134
rect 202726 236898 202768 237134
rect 202448 236866 202768 236898
rect 202448 201454 202768 201486
rect 202448 201218 202490 201454
rect 202726 201218 202768 201454
rect 202448 201134 202768 201218
rect 202448 200898 202490 201134
rect 202726 200898 202768 201134
rect 202448 200866 202768 200898
rect 202448 165454 202768 165486
rect 202448 165218 202490 165454
rect 202726 165218 202768 165454
rect 202448 165134 202768 165218
rect 202448 164898 202490 165134
rect 202726 164898 202768 165134
rect 202448 164866 202768 164898
rect 202448 129454 202768 129486
rect 202448 129218 202490 129454
rect 202726 129218 202768 129454
rect 202448 129134 202768 129218
rect 202448 128898 202490 129134
rect 202726 128898 202768 129134
rect 202448 128866 202768 128898
rect 202448 93454 202768 93486
rect 202448 93218 202490 93454
rect 202726 93218 202768 93454
rect 202448 93134 202768 93218
rect 202448 92898 202490 93134
rect 202726 92898 202768 93134
rect 202448 92866 202768 92898
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 197859 4180 197925 4181
rect 197859 4116 197860 4180
rect 197924 4116 197925 4180
rect 197859 4115 197925 4116
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 208902 13157 208962 542403
rect 210954 542000 211574 572058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 219203 699820 219269 699821
rect 219203 699756 219204 699820
rect 219268 699756 219269 699820
rect 219203 699755 219269 699756
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 542000 218414 542898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 217808 471454 218128 471486
rect 217808 471218 217850 471454
rect 218086 471218 218128 471454
rect 217808 471134 218128 471218
rect 217808 470898 217850 471134
rect 218086 470898 218128 471134
rect 217808 470866 218128 470898
rect 217808 435454 218128 435486
rect 217808 435218 217850 435454
rect 218086 435218 218128 435454
rect 217808 435134 218128 435218
rect 217808 434898 217850 435134
rect 218086 434898 218128 435134
rect 217808 434866 218128 434898
rect 217808 399454 218128 399486
rect 217808 399218 217850 399454
rect 218086 399218 218128 399454
rect 217808 399134 218128 399218
rect 217808 398898 217850 399134
rect 218086 398898 218128 399134
rect 217808 398866 218128 398898
rect 217808 363454 218128 363486
rect 217808 363218 217850 363454
rect 218086 363218 218128 363454
rect 217808 363134 218128 363218
rect 217808 362898 217850 363134
rect 218086 362898 218128 363134
rect 217808 362866 218128 362898
rect 217808 327454 218128 327486
rect 217808 327218 217850 327454
rect 218086 327218 218128 327454
rect 217808 327134 218128 327218
rect 217808 326898 217850 327134
rect 218086 326898 218128 327134
rect 217808 326866 218128 326898
rect 211294 301018 211354 303502
rect 217808 291454 218128 291486
rect 217808 291218 217850 291454
rect 218086 291218 218128 291454
rect 217808 291134 218128 291218
rect 217808 290898 217850 291134
rect 218086 290898 218128 291134
rect 217808 290866 218128 290898
rect 217808 255454 218128 255486
rect 217808 255218 217850 255454
rect 218086 255218 218128 255454
rect 217808 255134 218128 255218
rect 217808 254898 217850 255134
rect 218086 254898 218128 255134
rect 217808 254866 218128 254898
rect 217808 219454 218128 219486
rect 217808 219218 217850 219454
rect 218086 219218 218128 219454
rect 217808 219134 218128 219218
rect 217808 218898 217850 219134
rect 218086 218898 218128 219134
rect 217808 218866 218128 218898
rect 217808 183454 218128 183486
rect 217808 183218 217850 183454
rect 218086 183218 218128 183454
rect 217808 183134 218128 183218
rect 217808 182898 217850 183134
rect 218086 182898 218128 183134
rect 217808 182866 218128 182898
rect 217808 147454 218128 147486
rect 217808 147218 217850 147454
rect 218086 147218 218128 147454
rect 217808 147134 218128 147218
rect 217808 146898 217850 147134
rect 218086 146898 218128 147134
rect 217808 146866 218128 146898
rect 217808 111454 218128 111486
rect 217808 111218 217850 111454
rect 218086 111218 218128 111454
rect 217808 111134 218128 111218
rect 217808 110898 217850 111134
rect 218086 110898 218128 111134
rect 217808 110866 218128 110898
rect 217808 75454 218128 75486
rect 217808 75218 217850 75454
rect 218086 75218 218128 75454
rect 217808 75134 218128 75218
rect 217808 74898 217850 75134
rect 218086 74898 218128 75134
rect 217808 74866 218128 74898
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 208899 13156 208965 13157
rect 208899 13092 208900 13156
rect 208964 13092 208965 13156
rect 208899 13091 208965 13092
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 219206 57901 219266 699755
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 542000 222134 546618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 222699 542604 222765 542605
rect 222699 542540 222700 542604
rect 222764 542540 222765 542604
rect 222699 542539 222765 542540
rect 219939 539612 220005 539613
rect 219939 539548 219940 539612
rect 220004 539548 220005 539612
rect 219939 539547 220005 539548
rect 219203 57900 219269 57901
rect 219203 57836 219204 57900
rect 219268 57836 219269 57900
rect 219203 57835 219269 57836
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 219942 24173 220002 539547
rect 220310 301018 220370 303502
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 219939 24172 220005 24173
rect 219939 24108 219940 24172
rect 220004 24108 220005 24172
rect 219939 24107 220005 24108
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 42618
rect 222702 15877 222762 542539
rect 225234 542000 225854 550338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228219 543284 228285 543285
rect 228219 543220 228220 543284
rect 228284 543220 228285 543284
rect 228219 543219 228285 543220
rect 223619 539476 223685 539477
rect 223619 539412 223620 539476
rect 223684 539412 223685 539476
rect 223619 539411 223685 539412
rect 222699 15876 222765 15877
rect 222699 15812 222700 15876
rect 222764 15812 222765 15876
rect 222699 15811 222765 15812
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 223622 2957 223682 539411
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 228222 11797 228282 543219
rect 228954 542000 229574 554058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 230979 543148 231045 543149
rect 230979 543084 230980 543148
rect 231044 543084 231045 543148
rect 230979 543083 231045 543084
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228219 11796 228285 11797
rect 228219 11732 228220 11796
rect 228284 11732 228285 11796
rect 228219 11731 228285 11732
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 223619 2956 223685 2957
rect 223619 2892 223620 2956
rect 223684 2892 223685 2956
rect 223619 2891 223685 2892
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 230982 4181 231042 543083
rect 235794 542000 236414 560898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 237971 542468 238037 542469
rect 237971 542404 237972 542468
rect 238036 542404 238037 542468
rect 237971 542403 238037 542404
rect 233168 525454 233488 525486
rect 233168 525218 233210 525454
rect 233446 525218 233488 525454
rect 233168 525134 233488 525218
rect 233168 524898 233210 525134
rect 233446 524898 233488 525134
rect 233168 524866 233488 524898
rect 233168 489454 233488 489486
rect 233168 489218 233210 489454
rect 233446 489218 233488 489454
rect 233168 489134 233488 489218
rect 233168 488898 233210 489134
rect 233446 488898 233488 489134
rect 233168 488866 233488 488898
rect 233168 453454 233488 453486
rect 233168 453218 233210 453454
rect 233446 453218 233488 453454
rect 233168 453134 233488 453218
rect 233168 452898 233210 453134
rect 233446 452898 233488 453134
rect 233168 452866 233488 452898
rect 233168 417454 233488 417486
rect 233168 417218 233210 417454
rect 233446 417218 233488 417454
rect 233168 417134 233488 417218
rect 233168 416898 233210 417134
rect 233446 416898 233488 417134
rect 233168 416866 233488 416898
rect 233168 381454 233488 381486
rect 233168 381218 233210 381454
rect 233446 381218 233488 381454
rect 233168 381134 233488 381218
rect 233168 380898 233210 381134
rect 233446 380898 233488 381134
rect 233168 380866 233488 380898
rect 233168 345454 233488 345486
rect 233168 345218 233210 345454
rect 233446 345218 233488 345454
rect 233168 345134 233488 345218
rect 233168 344898 233210 345134
rect 233446 344898 233488 345134
rect 233168 344866 233488 344898
rect 233168 309454 233488 309486
rect 233168 309218 233210 309454
rect 233446 309218 233488 309454
rect 233168 309134 233488 309218
rect 233168 308898 233210 309134
rect 233446 308898 233488 309134
rect 233168 308866 233488 308898
rect 233168 273454 233488 273486
rect 233168 273218 233210 273454
rect 233446 273218 233488 273454
rect 233168 273134 233488 273218
rect 233168 272898 233210 273134
rect 233446 272898 233488 273134
rect 233168 272866 233488 272898
rect 233168 237454 233488 237486
rect 233168 237218 233210 237454
rect 233446 237218 233488 237454
rect 233168 237134 233488 237218
rect 233168 236898 233210 237134
rect 233446 236898 233488 237134
rect 233168 236866 233488 236898
rect 233168 201454 233488 201486
rect 233168 201218 233210 201454
rect 233446 201218 233488 201454
rect 233168 201134 233488 201218
rect 233168 200898 233210 201134
rect 233446 200898 233488 201134
rect 233168 200866 233488 200898
rect 233168 165454 233488 165486
rect 233168 165218 233210 165454
rect 233446 165218 233488 165454
rect 233168 165134 233488 165218
rect 233168 164898 233210 165134
rect 233446 164898 233488 165134
rect 233168 164866 233488 164898
rect 233168 129454 233488 129486
rect 233168 129218 233210 129454
rect 233446 129218 233488 129454
rect 233168 129134 233488 129218
rect 233168 128898 233210 129134
rect 233446 128898 233488 129134
rect 233168 128866 233488 128898
rect 233168 93454 233488 93486
rect 233168 93218 233210 93454
rect 233446 93218 233488 93454
rect 233168 93134 233488 93218
rect 233168 92898 233210 93134
rect 233446 92898 233488 93134
rect 233168 92866 233488 92898
rect 235794 57454 236414 58000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 230979 4180 231045 4181
rect 230979 4116 230980 4180
rect 231044 4116 231045 4180
rect 230979 4115 231045 4116
rect 235794 -1306 236414 20898
rect 237974 11797 238034 542403
rect 239514 542000 240134 564618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 242019 542604 242085 542605
rect 242019 542540 242020 542604
rect 242084 542540 242085 542604
rect 242019 542539 242085 542540
rect 240363 539476 240429 539477
rect 240363 539412 240364 539476
rect 240428 539412 240429 539476
rect 240363 539411 240429 539412
rect 239514 25174 240134 58000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 237971 11796 238037 11797
rect 237971 11732 237972 11796
rect 238036 11732 238037 11796
rect 237971 11731 238037 11732
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 -3226 240134 24618
rect 240366 17509 240426 539411
rect 240363 17508 240429 17509
rect 240363 17444 240364 17508
rect 240428 17444 240429 17508
rect 240363 17443 240429 17444
rect 242022 12069 242082 542539
rect 243234 542000 243854 568338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 542000 247574 572058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 251771 543692 251837 543693
rect 251771 543628 251772 543692
rect 251836 543628 251837 543692
rect 251771 543627 251837 543628
rect 250299 542468 250365 542469
rect 250299 542404 250300 542468
rect 250364 542404 250365 542468
rect 250299 542403 250365 542404
rect 246251 539612 246317 539613
rect 246251 539548 246252 539612
rect 246316 539548 246317 539612
rect 246251 539547 246317 539548
rect 243234 28894 243854 58000
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 242019 12068 242085 12069
rect 242019 12004 242020 12068
rect 242084 12004 242085 12068
rect 242019 12003 242085 12004
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28338
rect 246254 10301 246314 539547
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 248528 471454 248848 471486
rect 248528 471218 248570 471454
rect 248806 471218 248848 471454
rect 248528 471134 248848 471218
rect 248528 470898 248570 471134
rect 248806 470898 248848 471134
rect 248528 470866 248848 470898
rect 248528 435454 248848 435486
rect 248528 435218 248570 435454
rect 248806 435218 248848 435454
rect 248528 435134 248848 435218
rect 248528 434898 248570 435134
rect 248806 434898 248848 435134
rect 248528 434866 248848 434898
rect 248528 399454 248848 399486
rect 248528 399218 248570 399454
rect 248806 399218 248848 399454
rect 248528 399134 248848 399218
rect 248528 398898 248570 399134
rect 248806 398898 248848 399134
rect 248528 398866 248848 398898
rect 248528 363454 248848 363486
rect 248528 363218 248570 363454
rect 248806 363218 248848 363454
rect 248528 363134 248848 363218
rect 248528 362898 248570 363134
rect 248806 362898 248848 363134
rect 248528 362866 248848 362898
rect 248528 327454 248848 327486
rect 248528 327218 248570 327454
rect 248806 327218 248848 327454
rect 248528 327134 248848 327218
rect 248528 326898 248570 327134
rect 248806 326898 248848 327134
rect 248528 326866 248848 326898
rect 249382 301018 249442 303502
rect 248528 291454 248848 291486
rect 248528 291218 248570 291454
rect 248806 291218 248848 291454
rect 248528 291134 248848 291218
rect 248528 290898 248570 291134
rect 248806 290898 248848 291134
rect 248528 290866 248848 290898
rect 248528 255454 248848 255486
rect 248528 255218 248570 255454
rect 248806 255218 248848 255454
rect 248528 255134 248848 255218
rect 248528 254898 248570 255134
rect 248806 254898 248848 255134
rect 248528 254866 248848 254898
rect 248528 219454 248848 219486
rect 248528 219218 248570 219454
rect 248806 219218 248848 219454
rect 248528 219134 248848 219218
rect 248528 218898 248570 219134
rect 248806 218898 248848 219134
rect 248528 218866 248848 218898
rect 248528 183454 248848 183486
rect 248528 183218 248570 183454
rect 248806 183218 248848 183454
rect 248528 183134 248848 183218
rect 248528 182898 248570 183134
rect 248806 182898 248848 183134
rect 248528 182866 248848 182898
rect 248528 147454 248848 147486
rect 248528 147218 248570 147454
rect 248806 147218 248848 147454
rect 248528 147134 248848 147218
rect 248528 146898 248570 147134
rect 248806 146898 248848 147134
rect 248528 146866 248848 146898
rect 248528 111454 248848 111486
rect 248528 111218 248570 111454
rect 248806 111218 248848 111454
rect 248528 111134 248848 111218
rect 248528 110898 248570 111134
rect 248806 110898 248848 111134
rect 248528 110866 248848 110898
rect 248528 75454 248848 75486
rect 248528 75218 248570 75454
rect 248806 75218 248848 75454
rect 248528 75134 248848 75218
rect 248528 74898 248570 75134
rect 248806 74898 248848 75134
rect 248528 74866 248848 74898
rect 246954 32614 247574 58000
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 246251 10300 246317 10301
rect 246251 10236 246252 10300
rect 246316 10236 246317 10300
rect 246251 10235 246317 10236
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 250302 5677 250362 542403
rect 251774 21317 251834 543627
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 255819 543148 255885 543149
rect 255819 543084 255820 543148
rect 255884 543084 255885 543148
rect 255819 543083 255885 543084
rect 253794 542000 254414 542898
rect 252507 539612 252573 539613
rect 252507 539548 252508 539612
rect 252572 539548 252573 539612
rect 252507 539547 252573 539548
rect 251771 21316 251837 21317
rect 251771 21252 251772 21316
rect 251836 21252 251837 21316
rect 251771 21251 251837 21252
rect 250299 5676 250365 5677
rect 250299 5612 250300 5676
rect 250364 5612 250365 5676
rect 250299 5611 250365 5612
rect 252510 3229 252570 539547
rect 253794 39454 254414 58000
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 255822 10981 255882 543083
rect 257514 542000 258134 546618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 542000 261854 550338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 542000 265574 554058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271091 542876 271157 542877
rect 271091 542812 271092 542876
rect 271156 542812 271157 542876
rect 271091 542811 271157 542812
rect 266859 542604 266925 542605
rect 266859 542540 266860 542604
rect 266924 542540 266925 542604
rect 266859 542539 266925 542540
rect 263888 525454 264208 525486
rect 263888 525218 263930 525454
rect 264166 525218 264208 525454
rect 263888 525134 264208 525218
rect 263888 524898 263930 525134
rect 264166 524898 264208 525134
rect 263888 524866 264208 524898
rect 263888 489454 264208 489486
rect 263888 489218 263930 489454
rect 264166 489218 264208 489454
rect 263888 489134 264208 489218
rect 263888 488898 263930 489134
rect 264166 488898 264208 489134
rect 263888 488866 264208 488898
rect 263888 453454 264208 453486
rect 263888 453218 263930 453454
rect 264166 453218 264208 453454
rect 263888 453134 264208 453218
rect 263888 452898 263930 453134
rect 264166 452898 264208 453134
rect 263888 452866 264208 452898
rect 263888 417454 264208 417486
rect 263888 417218 263930 417454
rect 264166 417218 264208 417454
rect 263888 417134 264208 417218
rect 263888 416898 263930 417134
rect 264166 416898 264208 417134
rect 263888 416866 264208 416898
rect 263888 381454 264208 381486
rect 263888 381218 263930 381454
rect 264166 381218 264208 381454
rect 263888 381134 264208 381218
rect 263888 380898 263930 381134
rect 264166 380898 264208 381134
rect 263888 380866 264208 380898
rect 263888 345454 264208 345486
rect 263888 345218 263930 345454
rect 264166 345218 264208 345454
rect 263888 345134 264208 345218
rect 263888 344898 263930 345134
rect 264166 344898 264208 345134
rect 263888 344866 264208 344898
rect 263888 309454 264208 309486
rect 263888 309218 263930 309454
rect 264166 309218 264208 309454
rect 263888 309134 264208 309218
rect 263888 308898 263930 309134
rect 264166 308898 264208 309134
rect 263888 308866 264208 308898
rect 263888 273454 264208 273486
rect 263888 273218 263930 273454
rect 264166 273218 264208 273454
rect 263888 273134 264208 273218
rect 263888 272898 263930 273134
rect 264166 272898 264208 273134
rect 263888 272866 264208 272898
rect 263888 237454 264208 237486
rect 263888 237218 263930 237454
rect 264166 237218 264208 237454
rect 263888 237134 264208 237218
rect 263888 236898 263930 237134
rect 264166 236898 264208 237134
rect 263888 236866 264208 236898
rect 263888 201454 264208 201486
rect 263888 201218 263930 201454
rect 264166 201218 264208 201454
rect 263888 201134 264208 201218
rect 263888 200898 263930 201134
rect 264166 200898 264208 201134
rect 263888 200866 264208 200898
rect 263888 165454 264208 165486
rect 263888 165218 263930 165454
rect 264166 165218 264208 165454
rect 263888 165134 264208 165218
rect 263888 164898 263930 165134
rect 264166 164898 264208 165134
rect 263888 164866 264208 164898
rect 263888 129454 264208 129486
rect 263888 129218 263930 129454
rect 264166 129218 264208 129454
rect 263888 129134 264208 129218
rect 263888 128898 263930 129134
rect 264166 128898 264208 129134
rect 263888 128866 264208 128898
rect 263888 93454 264208 93486
rect 263888 93218 263930 93454
rect 264166 93218 264208 93454
rect 263888 93134 264208 93218
rect 263888 92898 263930 93134
rect 264166 92898 264208 93134
rect 263888 92866 264208 92898
rect 257514 43174 258134 58000
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 255819 10980 255885 10981
rect 255819 10916 255820 10980
rect 255884 10916 255885 10980
rect 255819 10915 255885 10916
rect 252507 3228 252573 3229
rect 252507 3164 252508 3228
rect 252572 3164 252573 3228
rect 252507 3163 252573 3164
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 266862 5677 266922 542539
rect 269619 539476 269685 539477
rect 269619 539412 269620 539476
rect 269684 539412 269685 539476
rect 269619 539411 269685 539412
rect 267966 301018 268026 303502
rect 269622 21453 269682 539411
rect 269619 21452 269685 21453
rect 269619 21388 269620 21452
rect 269684 21388 269685 21452
rect 269619 21387 269685 21388
rect 266859 5676 266925 5677
rect 266859 5612 266860 5676
rect 266924 5612 266925 5676
rect 266859 5611 266925 5612
rect 271094 4181 271154 542811
rect 271794 542000 272414 560898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 542000 276134 564618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 277899 543556 277965 543557
rect 277899 543492 277900 543556
rect 277964 543492 277965 543556
rect 277899 543491 277965 543492
rect 271794 57454 272414 58000
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271091 4180 271157 4181
rect 271091 4116 271092 4180
rect 271156 4116 271157 4180
rect 271091 4115 271157 4116
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 277902 4181 277962 543491
rect 279234 542000 279854 568338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 280659 543012 280725 543013
rect 280659 542948 280660 543012
rect 280724 542948 280725 543012
rect 280659 542947 280725 542948
rect 279003 539476 279069 539477
rect 279003 539412 279004 539476
rect 279068 539412 279069 539476
rect 279003 539411 279069 539412
rect 277899 4180 277965 4181
rect 277899 4116 277900 4180
rect 277964 4116 277965 4180
rect 277899 4115 277965 4116
rect 279006 3229 279066 539411
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 279248 471454 279568 471486
rect 279248 471218 279290 471454
rect 279526 471218 279568 471454
rect 279248 471134 279568 471218
rect 279248 470898 279290 471134
rect 279526 470898 279568 471134
rect 279248 470866 279568 470898
rect 279248 435454 279568 435486
rect 279248 435218 279290 435454
rect 279526 435218 279568 435454
rect 279248 435134 279568 435218
rect 279248 434898 279290 435134
rect 279526 434898 279568 435134
rect 279248 434866 279568 434898
rect 279248 399454 279568 399486
rect 279248 399218 279290 399454
rect 279526 399218 279568 399454
rect 279248 399134 279568 399218
rect 279248 398898 279290 399134
rect 279526 398898 279568 399134
rect 279248 398866 279568 398898
rect 279248 363454 279568 363486
rect 279248 363218 279290 363454
rect 279526 363218 279568 363454
rect 279248 363134 279568 363218
rect 279248 362898 279290 363134
rect 279526 362898 279568 363134
rect 279248 362866 279568 362898
rect 279248 327454 279568 327486
rect 279248 327218 279290 327454
rect 279526 327218 279568 327454
rect 279248 327134 279568 327218
rect 279248 326898 279290 327134
rect 279526 326898 279568 327134
rect 279248 326866 279568 326898
rect 279248 291454 279568 291486
rect 279248 291218 279290 291454
rect 279526 291218 279568 291454
rect 279248 291134 279568 291218
rect 279248 290898 279290 291134
rect 279526 290898 279568 291134
rect 279248 290866 279568 290898
rect 279248 255454 279568 255486
rect 279248 255218 279290 255454
rect 279526 255218 279568 255454
rect 279248 255134 279568 255218
rect 279248 254898 279290 255134
rect 279526 254898 279568 255134
rect 279248 254866 279568 254898
rect 279248 219454 279568 219486
rect 279248 219218 279290 219454
rect 279526 219218 279568 219454
rect 279248 219134 279568 219218
rect 279248 218898 279290 219134
rect 279526 218898 279568 219134
rect 279248 218866 279568 218898
rect 279248 183454 279568 183486
rect 279248 183218 279290 183454
rect 279526 183218 279568 183454
rect 279248 183134 279568 183218
rect 279248 182898 279290 183134
rect 279526 182898 279568 183134
rect 279248 182866 279568 182898
rect 279248 147454 279568 147486
rect 279248 147218 279290 147454
rect 279526 147218 279568 147454
rect 279248 147134 279568 147218
rect 279248 146898 279290 147134
rect 279526 146898 279568 147134
rect 279248 146866 279568 146898
rect 279248 111454 279568 111486
rect 279248 111218 279290 111454
rect 279526 111218 279568 111454
rect 279248 111134 279568 111218
rect 279248 110898 279290 111134
rect 279526 110898 279568 111134
rect 279248 110866 279568 110898
rect 279248 75454 279568 75486
rect 279248 75218 279290 75454
rect 279526 75218 279568 75454
rect 279248 75134 279568 75218
rect 279248 74898 279290 75134
rect 279526 74898 279568 75134
rect 279248 74866 279568 74898
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279003 3228 279069 3229
rect 279003 3164 279004 3228
rect 279068 3164 279069 3228
rect 279003 3163 279069 3164
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 28338
rect 280662 10437 280722 542947
rect 282954 542000 283574 572058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 542000 290414 542898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 542000 294134 546618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 542000 297854 550338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 542000 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 542000 308414 560898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 542000 312134 564618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 542000 315854 568338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 542000 319574 572058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 327579 543420 327645 543421
rect 327579 543356 327580 543420
rect 327644 543356 327645 543420
rect 327579 543355 327645 543356
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 322059 542876 322125 542877
rect 322059 542812 322060 542876
rect 322124 542812 322125 542876
rect 322059 542811 322125 542812
rect 304947 541108 305013 541109
rect 304947 541044 304948 541108
rect 305012 541044 305013 541108
rect 304947 541043 305013 541044
rect 283787 539612 283853 539613
rect 283787 539548 283788 539612
rect 283852 539548 283853 539612
rect 283787 539547 283853 539548
rect 282954 32614 283574 58000
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 280659 10436 280725 10437
rect 280659 10372 280660 10436
rect 280724 10372 280725 10436
rect 280659 10371 280725 10372
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 283790 3093 283850 539547
rect 298139 539476 298205 539477
rect 298139 539412 298140 539476
rect 298204 539412 298205 539476
rect 298139 539411 298205 539412
rect 294608 525454 294928 525486
rect 294608 525218 294650 525454
rect 294886 525218 294928 525454
rect 294608 525134 294928 525218
rect 294608 524898 294650 525134
rect 294886 524898 294928 525134
rect 294608 524866 294928 524898
rect 294608 489454 294928 489486
rect 294608 489218 294650 489454
rect 294886 489218 294928 489454
rect 294608 489134 294928 489218
rect 294608 488898 294650 489134
rect 294886 488898 294928 489134
rect 294608 488866 294928 488898
rect 294608 453454 294928 453486
rect 294608 453218 294650 453454
rect 294886 453218 294928 453454
rect 294608 453134 294928 453218
rect 294608 452898 294650 453134
rect 294886 452898 294928 453134
rect 294608 452866 294928 452898
rect 294608 417454 294928 417486
rect 294608 417218 294650 417454
rect 294886 417218 294928 417454
rect 294608 417134 294928 417218
rect 294608 416898 294650 417134
rect 294886 416898 294928 417134
rect 294608 416866 294928 416898
rect 294608 381454 294928 381486
rect 294608 381218 294650 381454
rect 294886 381218 294928 381454
rect 294608 381134 294928 381218
rect 294608 380898 294650 381134
rect 294886 380898 294928 381134
rect 294608 380866 294928 380898
rect 294608 345454 294928 345486
rect 294608 345218 294650 345454
rect 294886 345218 294928 345454
rect 294608 345134 294928 345218
rect 294608 344898 294650 345134
rect 294886 344898 294928 345134
rect 294608 344866 294928 344898
rect 294608 309454 294928 309486
rect 294608 309218 294650 309454
rect 294886 309218 294928 309454
rect 294608 309134 294928 309218
rect 294608 308898 294650 309134
rect 294886 308898 294928 309134
rect 294608 308866 294928 308898
rect 287654 301018 287714 303502
rect 294608 273454 294928 273486
rect 294608 273218 294650 273454
rect 294886 273218 294928 273454
rect 294608 273134 294928 273218
rect 294608 272898 294650 273134
rect 294886 272898 294928 273134
rect 294608 272866 294928 272898
rect 294608 237454 294928 237486
rect 294608 237218 294650 237454
rect 294886 237218 294928 237454
rect 294608 237134 294928 237218
rect 294608 236898 294650 237134
rect 294886 236898 294928 237134
rect 294608 236866 294928 236898
rect 294608 201454 294928 201486
rect 294608 201218 294650 201454
rect 294886 201218 294928 201454
rect 294608 201134 294928 201218
rect 294608 200898 294650 201134
rect 294886 200898 294928 201134
rect 294608 200866 294928 200898
rect 294608 165454 294928 165486
rect 294608 165218 294650 165454
rect 294886 165218 294928 165454
rect 294608 165134 294928 165218
rect 294608 164898 294650 165134
rect 294886 164898 294928 165134
rect 294608 164866 294928 164898
rect 294608 129454 294928 129486
rect 294608 129218 294650 129454
rect 294886 129218 294928 129454
rect 294608 129134 294928 129218
rect 294608 128898 294650 129134
rect 294886 128898 294928 129134
rect 294608 128866 294928 128898
rect 294608 93454 294928 93486
rect 294608 93218 294650 93454
rect 294886 93218 294928 93454
rect 294608 93134 294928 93218
rect 294608 92898 294650 93134
rect 294886 92898 294928 93134
rect 294608 92866 294928 92898
rect 289794 39454 290414 58000
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 283787 3092 283853 3093
rect 283787 3028 283788 3092
rect 283852 3028 283853 3092
rect 283787 3027 283853 3028
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 298142 4045 298202 539411
rect 300954 50614 301574 58000
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 298139 4044 298205 4045
rect 298139 3980 298140 4044
rect 298204 3980 298205 4044
rect 298139 3979 298205 3980
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 304950 3093 305010 541043
rect 313227 539612 313293 539613
rect 313227 539548 313228 539612
rect 313292 539548 313293 539612
rect 313227 539547 313293 539548
rect 309179 539476 309245 539477
rect 309179 539412 309180 539476
rect 309244 539412 309245 539476
rect 309179 539411 309245 539412
rect 309182 325710 309242 539411
rect 309968 507454 310288 507486
rect 309968 507218 310010 507454
rect 310246 507218 310288 507454
rect 309968 507134 310288 507218
rect 309968 506898 310010 507134
rect 310246 506898 310288 507134
rect 309968 506866 310288 506898
rect 309968 471454 310288 471486
rect 309968 471218 310010 471454
rect 310246 471218 310288 471454
rect 309968 471134 310288 471218
rect 309968 470898 310010 471134
rect 310246 470898 310288 471134
rect 309968 470866 310288 470898
rect 309968 435454 310288 435486
rect 309968 435218 310010 435454
rect 310246 435218 310288 435454
rect 309968 435134 310288 435218
rect 309968 434898 310010 435134
rect 310246 434898 310288 435134
rect 309968 434866 310288 434898
rect 309968 399454 310288 399486
rect 309968 399218 310010 399454
rect 310246 399218 310288 399454
rect 309968 399134 310288 399218
rect 309968 398898 310010 399134
rect 310246 398898 310288 399134
rect 309968 398866 310288 398898
rect 309968 363454 310288 363486
rect 309968 363218 310010 363454
rect 310246 363218 310288 363454
rect 309968 363134 310288 363218
rect 309968 362898 310010 363134
rect 310246 362898 310288 363134
rect 309968 362866 310288 362898
rect 309968 327454 310288 327486
rect 309968 327218 310010 327454
rect 310246 327218 310288 327454
rect 309968 327134 310288 327218
rect 309968 326898 310010 327134
rect 310246 326898 310288 327134
rect 309968 326866 310288 326898
rect 309182 325650 309610 325710
rect 309550 296730 309610 325650
rect 309182 296670 309610 296730
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 304947 3092 305013 3093
rect 304947 3028 304948 3092
rect 305012 3028 305013 3092
rect 304947 3027 305013 3028
rect 307794 -1306 308414 20898
rect 309182 4538 309242 296670
rect 309968 291454 310288 291486
rect 309968 291218 310010 291454
rect 310246 291218 310288 291454
rect 309968 291134 310288 291218
rect 309968 290898 310010 291134
rect 310246 290898 310288 291134
rect 309968 290866 310288 290898
rect 309968 255454 310288 255486
rect 309968 255218 310010 255454
rect 310246 255218 310288 255454
rect 309968 255134 310288 255218
rect 309968 254898 310010 255134
rect 310246 254898 310288 255134
rect 309968 254866 310288 254898
rect 309968 219454 310288 219486
rect 309968 219218 310010 219454
rect 310246 219218 310288 219454
rect 309968 219134 310288 219218
rect 309968 218898 310010 219134
rect 310246 218898 310288 219134
rect 309968 218866 310288 218898
rect 309968 183454 310288 183486
rect 309968 183218 310010 183454
rect 310246 183218 310288 183454
rect 309968 183134 310288 183218
rect 309968 182898 310010 183134
rect 310246 182898 310288 183134
rect 309968 182866 310288 182898
rect 309968 147454 310288 147486
rect 309968 147218 310010 147454
rect 310246 147218 310288 147454
rect 309968 147134 310288 147218
rect 309968 146898 310010 147134
rect 310246 146898 310288 147134
rect 309968 146866 310288 146898
rect 309968 111454 310288 111486
rect 309968 111218 310010 111454
rect 310246 111218 310288 111454
rect 309968 111134 310288 111218
rect 309968 110898 310010 111134
rect 310246 110898 310288 111134
rect 309968 110866 310288 110898
rect 309968 75454 310288 75486
rect 309968 75218 310010 75454
rect 310246 75218 310288 75454
rect 309968 75134 310288 75218
rect 309968 74898 310010 75134
rect 310246 74898 310288 75134
rect 309968 74866 310288 74898
rect 311514 25174 312134 58000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 -3226 312134 24618
rect 313230 15877 313290 539547
rect 316542 301018 316602 303502
rect 315234 28894 315854 58000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 313227 15876 313293 15877
rect 313227 15812 313228 15876
rect 313292 15812 313293 15876
rect 313227 15811 313293 15812
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 322062 11661 322122 542811
rect 325794 542000 326414 542898
rect 325328 525454 325648 525486
rect 325328 525218 325370 525454
rect 325606 525218 325648 525454
rect 325328 525134 325648 525218
rect 325328 524898 325370 525134
rect 325606 524898 325648 525134
rect 325328 524866 325648 524898
rect 325328 489454 325648 489486
rect 325328 489218 325370 489454
rect 325606 489218 325648 489454
rect 325328 489134 325648 489218
rect 325328 488898 325370 489134
rect 325606 488898 325648 489134
rect 325328 488866 325648 488898
rect 325328 453454 325648 453486
rect 325328 453218 325370 453454
rect 325606 453218 325648 453454
rect 325328 453134 325648 453218
rect 325328 452898 325370 453134
rect 325606 452898 325648 453134
rect 325328 452866 325648 452898
rect 325328 417454 325648 417486
rect 325328 417218 325370 417454
rect 325606 417218 325648 417454
rect 325328 417134 325648 417218
rect 325328 416898 325370 417134
rect 325606 416898 325648 417134
rect 325328 416866 325648 416898
rect 325328 381454 325648 381486
rect 325328 381218 325370 381454
rect 325606 381218 325648 381454
rect 325328 381134 325648 381218
rect 325328 380898 325370 381134
rect 325606 380898 325648 381134
rect 325328 380866 325648 380898
rect 325328 345454 325648 345486
rect 325328 345218 325370 345454
rect 325606 345218 325648 345454
rect 325328 345134 325648 345218
rect 325328 344898 325370 345134
rect 325606 344898 325648 345134
rect 325328 344866 325648 344898
rect 325328 309454 325648 309486
rect 325328 309218 325370 309454
rect 325606 309218 325648 309454
rect 325328 309134 325648 309218
rect 325328 308898 325370 309134
rect 325606 308898 325648 309134
rect 325328 308866 325648 308898
rect 325328 273454 325648 273486
rect 325328 273218 325370 273454
rect 325606 273218 325648 273454
rect 325328 273134 325648 273218
rect 325328 272898 325370 273134
rect 325606 272898 325648 273134
rect 325328 272866 325648 272898
rect 325328 237454 325648 237486
rect 325328 237218 325370 237454
rect 325606 237218 325648 237454
rect 325328 237134 325648 237218
rect 325328 236898 325370 237134
rect 325606 236898 325648 237134
rect 325328 236866 325648 236898
rect 325328 201454 325648 201486
rect 325328 201218 325370 201454
rect 325606 201218 325648 201454
rect 325328 201134 325648 201218
rect 325328 200898 325370 201134
rect 325606 200898 325648 201134
rect 325328 200866 325648 200898
rect 325328 165454 325648 165486
rect 325328 165218 325370 165454
rect 325606 165218 325648 165454
rect 325328 165134 325648 165218
rect 325328 164898 325370 165134
rect 325606 164898 325648 165134
rect 325328 164866 325648 164898
rect 325328 129454 325648 129486
rect 325328 129218 325370 129454
rect 325606 129218 325648 129454
rect 325328 129134 325648 129218
rect 325328 128898 325370 129134
rect 325606 128898 325648 129134
rect 325328 128866 325648 128898
rect 325328 93454 325648 93486
rect 325328 93218 325370 93454
rect 325606 93218 325648 93454
rect 325328 93134 325648 93218
rect 325328 92898 325370 93134
rect 325606 92898 325648 93134
rect 325328 92866 325648 92898
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 322059 11660 322125 11661
rect 322059 11596 322060 11660
rect 322124 11596 322125 11660
rect 322059 11595 322125 11596
rect 325794 3454 326414 38898
rect 327582 10437 327642 543355
rect 329514 542000 330134 546618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 331811 543012 331877 543013
rect 331811 542948 331812 543012
rect 331876 542948 331877 543012
rect 331811 542947 331877 542948
rect 330339 539612 330405 539613
rect 330339 539548 330340 539612
rect 330404 539548 330405 539612
rect 330339 539547 330405 539548
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 327579 10436 327645 10437
rect 327579 10372 327580 10436
rect 327644 10372 327645 10436
rect 327579 10371 327645 10372
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 330342 3093 330402 539547
rect 331814 4181 331874 542947
rect 333234 542000 333854 550338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 335859 543012 335925 543013
rect 335859 542948 335860 543012
rect 335924 542948 335925 543012
rect 335859 542947 335925 542948
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 331811 4180 331877 4181
rect 331811 4116 331812 4180
rect 331876 4116 331877 4180
rect 331811 4115 331877 4116
rect 330339 3092 330405 3093
rect 330339 3028 330340 3092
rect 330404 3028 330405 3092
rect 330339 3027 330405 3028
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 10338
rect 335862 5677 335922 542947
rect 336954 542000 337574 554058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 542000 344414 560898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 542000 348134 564618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 542000 351854 568338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 353891 542604 353957 542605
rect 353891 542540 353892 542604
rect 353956 542540 353957 542604
rect 353891 542539 353957 542540
rect 341195 539612 341261 539613
rect 341195 539548 341196 539612
rect 341260 539548 341261 539612
rect 341195 539547 341261 539548
rect 340688 507454 341008 507486
rect 340688 507218 340730 507454
rect 340966 507218 341008 507454
rect 340688 507134 341008 507218
rect 340688 506898 340730 507134
rect 340966 506898 341008 507134
rect 340688 506866 341008 506898
rect 340688 471454 341008 471486
rect 340688 471218 340730 471454
rect 340966 471218 341008 471454
rect 340688 471134 341008 471218
rect 340688 470898 340730 471134
rect 340966 470898 341008 471134
rect 340688 470866 341008 470898
rect 340688 435454 341008 435486
rect 340688 435218 340730 435454
rect 340966 435218 341008 435454
rect 340688 435134 341008 435218
rect 340688 434898 340730 435134
rect 340966 434898 341008 435134
rect 340688 434866 341008 434898
rect 340688 399454 341008 399486
rect 340688 399218 340730 399454
rect 340966 399218 341008 399454
rect 340688 399134 341008 399218
rect 340688 398898 340730 399134
rect 340966 398898 341008 399134
rect 340688 398866 341008 398898
rect 340688 363454 341008 363486
rect 340688 363218 340730 363454
rect 340966 363218 341008 363454
rect 340688 363134 341008 363218
rect 340688 362898 340730 363134
rect 340966 362898 341008 363134
rect 340688 362866 341008 362898
rect 340688 327454 341008 327486
rect 340688 327218 340730 327454
rect 340966 327218 341008 327454
rect 340688 327134 341008 327218
rect 340688 326898 340730 327134
rect 340966 326898 341008 327134
rect 340688 326866 341008 326898
rect 340688 291454 341008 291486
rect 340688 291218 340730 291454
rect 340966 291218 341008 291454
rect 340688 291134 341008 291218
rect 340688 290898 340730 291134
rect 340966 290898 341008 291134
rect 340688 290866 341008 290898
rect 340688 255454 341008 255486
rect 340688 255218 340730 255454
rect 340966 255218 341008 255454
rect 340688 255134 341008 255218
rect 340688 254898 340730 255134
rect 340966 254898 341008 255134
rect 340688 254866 341008 254898
rect 340688 219454 341008 219486
rect 340688 219218 340730 219454
rect 340966 219218 341008 219454
rect 340688 219134 341008 219218
rect 340688 218898 340730 219134
rect 340966 218898 341008 219134
rect 340688 218866 341008 218898
rect 340688 183454 341008 183486
rect 340688 183218 340730 183454
rect 340966 183218 341008 183454
rect 340688 183134 341008 183218
rect 340688 182898 340730 183134
rect 340966 182898 341008 183134
rect 340688 182866 341008 182898
rect 340688 147454 341008 147486
rect 340688 147218 340730 147454
rect 340966 147218 341008 147454
rect 340688 147134 341008 147218
rect 340688 146898 340730 147134
rect 340966 146898 341008 147134
rect 340688 146866 341008 146898
rect 340688 111454 341008 111486
rect 340688 111218 340730 111454
rect 340966 111218 341008 111454
rect 340688 111134 341008 111218
rect 340688 110898 340730 111134
rect 340966 110898 341008 111134
rect 340688 110866 341008 110898
rect 340688 75454 341008 75486
rect 340688 75218 340730 75454
rect 340966 75218 341008 75454
rect 340688 75134 341008 75218
rect 340688 74898 340730 75134
rect 340966 74898 341008 75134
rect 340688 74866 341008 74898
rect 336954 50614 337574 58000
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 335859 5676 335925 5677
rect 335859 5612 335860 5676
rect 335924 5612 335925 5676
rect 335859 5611 335925 5612
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 341198 9621 341258 539547
rect 350395 539476 350461 539477
rect 350395 539412 350396 539476
rect 350460 539412 350461 539476
rect 350395 539411 350461 539412
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 341195 9620 341261 9621
rect 341195 9556 341196 9620
rect 341260 9556 341261 9620
rect 341195 9555 341261 9556
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 350398 3093 350458 539411
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 350395 3092 350461 3093
rect 350395 3028 350396 3092
rect 350460 3028 350461 3092
rect 350395 3027 350461 3028
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 28338
rect 353894 15877 353954 542539
rect 354954 542000 355574 572058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 542000 362414 542898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 363459 542876 363525 542877
rect 363459 542812 363460 542876
rect 363524 542812 363525 542876
rect 363459 542811 363525 542812
rect 360699 539612 360765 539613
rect 360699 539548 360700 539612
rect 360764 539548 360765 539612
rect 360699 539547 360765 539548
rect 356048 525454 356368 525486
rect 356048 525218 356090 525454
rect 356326 525218 356368 525454
rect 356048 525134 356368 525218
rect 356048 524898 356090 525134
rect 356326 524898 356368 525134
rect 356048 524866 356368 524898
rect 356048 489454 356368 489486
rect 356048 489218 356090 489454
rect 356326 489218 356368 489454
rect 356048 489134 356368 489218
rect 356048 488898 356090 489134
rect 356326 488898 356368 489134
rect 356048 488866 356368 488898
rect 356048 453454 356368 453486
rect 356048 453218 356090 453454
rect 356326 453218 356368 453454
rect 356048 453134 356368 453218
rect 356048 452898 356090 453134
rect 356326 452898 356368 453134
rect 356048 452866 356368 452898
rect 356048 417454 356368 417486
rect 356048 417218 356090 417454
rect 356326 417218 356368 417454
rect 356048 417134 356368 417218
rect 356048 416898 356090 417134
rect 356326 416898 356368 417134
rect 356048 416866 356368 416898
rect 356048 381454 356368 381486
rect 356048 381218 356090 381454
rect 356326 381218 356368 381454
rect 356048 381134 356368 381218
rect 356048 380898 356090 381134
rect 356326 380898 356368 381134
rect 356048 380866 356368 380898
rect 356048 345454 356368 345486
rect 356048 345218 356090 345454
rect 356326 345218 356368 345454
rect 356048 345134 356368 345218
rect 356048 344898 356090 345134
rect 356326 344898 356368 345134
rect 356048 344866 356368 344898
rect 356048 309454 356368 309486
rect 356048 309218 356090 309454
rect 356326 309218 356368 309454
rect 356048 309134 356368 309218
rect 356048 308898 356090 309134
rect 356326 308898 356368 309134
rect 356048 308866 356368 308898
rect 354998 301018 355058 303502
rect 356048 273454 356368 273486
rect 356048 273218 356090 273454
rect 356326 273218 356368 273454
rect 356048 273134 356368 273218
rect 356048 272898 356090 273134
rect 356326 272898 356368 273134
rect 356048 272866 356368 272898
rect 356048 237454 356368 237486
rect 356048 237218 356090 237454
rect 356326 237218 356368 237454
rect 356048 237134 356368 237218
rect 356048 236898 356090 237134
rect 356326 236898 356368 237134
rect 356048 236866 356368 236898
rect 356048 201454 356368 201486
rect 356048 201218 356090 201454
rect 356326 201218 356368 201454
rect 356048 201134 356368 201218
rect 356048 200898 356090 201134
rect 356326 200898 356368 201134
rect 356048 200866 356368 200898
rect 356048 165454 356368 165486
rect 356048 165218 356090 165454
rect 356326 165218 356368 165454
rect 356048 165134 356368 165218
rect 356048 164898 356090 165134
rect 356326 164898 356368 165134
rect 356048 164866 356368 164898
rect 356048 129454 356368 129486
rect 356048 129218 356090 129454
rect 356326 129218 356368 129454
rect 356048 129134 356368 129218
rect 356048 128898 356090 129134
rect 356326 128898 356368 129134
rect 356048 128866 356368 128898
rect 356048 93454 356368 93486
rect 356048 93218 356090 93454
rect 356326 93218 356368 93454
rect 356048 93134 356368 93218
rect 356048 92898 356090 93134
rect 356326 92898 356368 93134
rect 356048 92866 356368 92898
rect 354954 32614 355574 58000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 353891 15876 353957 15877
rect 353891 15812 353892 15876
rect 353956 15812 353957 15876
rect 353891 15811 353957 15812
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 360702 2957 360762 539547
rect 361794 39454 362414 58000
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 363462 14653 363522 542811
rect 365514 542000 366134 546618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 367691 542740 367757 542741
rect 367691 542676 367692 542740
rect 367756 542676 367757 542740
rect 367691 542675 367757 542676
rect 365514 43174 366134 58000
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 363459 14652 363525 14653
rect 363459 14588 363460 14652
rect 363524 14588 363525 14652
rect 363459 14587 363525 14588
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 360699 2956 360765 2957
rect 360699 2892 360700 2956
rect 360764 2892 360765 2956
rect 360699 2891 360765 2892
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 42618
rect 367694 40629 367754 542675
rect 369234 542000 369854 550338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 542000 373574 554058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 542000 380414 560898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 542000 384134 564618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 542000 387854 568338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 389771 542604 389837 542605
rect 389771 542540 389772 542604
rect 389836 542540 389837 542604
rect 389771 542539 389837 542540
rect 377259 539612 377325 539613
rect 377259 539548 377260 539612
rect 377324 539548 377325 539612
rect 377259 539547 377325 539548
rect 382227 539612 382293 539613
rect 382227 539548 382228 539612
rect 382292 539548 382293 539612
rect 382227 539547 382293 539548
rect 384987 539612 385053 539613
rect 384987 539548 384988 539612
rect 385052 539548 385053 539612
rect 384987 539547 385053 539548
rect 387931 539612 387997 539613
rect 387931 539548 387932 539612
rect 387996 539548 387997 539612
rect 387931 539547 387997 539548
rect 371408 507454 371728 507486
rect 371408 507218 371450 507454
rect 371686 507218 371728 507454
rect 371408 507134 371728 507218
rect 371408 506898 371450 507134
rect 371686 506898 371728 507134
rect 371408 506866 371728 506898
rect 371408 471454 371728 471486
rect 371408 471218 371450 471454
rect 371686 471218 371728 471454
rect 371408 471134 371728 471218
rect 371408 470898 371450 471134
rect 371686 470898 371728 471134
rect 371408 470866 371728 470898
rect 371408 435454 371728 435486
rect 371408 435218 371450 435454
rect 371686 435218 371728 435454
rect 371408 435134 371728 435218
rect 371408 434898 371450 435134
rect 371686 434898 371728 435134
rect 371408 434866 371728 434898
rect 371408 399454 371728 399486
rect 371408 399218 371450 399454
rect 371686 399218 371728 399454
rect 371408 399134 371728 399218
rect 371408 398898 371450 399134
rect 371686 398898 371728 399134
rect 371408 398866 371728 398898
rect 371408 363454 371728 363486
rect 371408 363218 371450 363454
rect 371686 363218 371728 363454
rect 371408 363134 371728 363218
rect 371408 362898 371450 363134
rect 371686 362898 371728 363134
rect 371408 362866 371728 362898
rect 371408 327454 371728 327486
rect 371408 327218 371450 327454
rect 371686 327218 371728 327454
rect 371408 327134 371728 327218
rect 371408 326898 371450 327134
rect 371686 326898 371728 327134
rect 371408 326866 371728 326898
rect 374134 301018 374194 303502
rect 371408 291454 371728 291486
rect 371408 291218 371450 291454
rect 371686 291218 371728 291454
rect 371408 291134 371728 291218
rect 371408 290898 371450 291134
rect 371686 290898 371728 291134
rect 371408 290866 371728 290898
rect 371408 255454 371728 255486
rect 371408 255218 371450 255454
rect 371686 255218 371728 255454
rect 371408 255134 371728 255218
rect 371408 254898 371450 255134
rect 371686 254898 371728 255134
rect 371408 254866 371728 254898
rect 371408 219454 371728 219486
rect 371408 219218 371450 219454
rect 371686 219218 371728 219454
rect 371408 219134 371728 219218
rect 371408 218898 371450 219134
rect 371686 218898 371728 219134
rect 371408 218866 371728 218898
rect 371408 183454 371728 183486
rect 371408 183218 371450 183454
rect 371686 183218 371728 183454
rect 371408 183134 371728 183218
rect 371408 182898 371450 183134
rect 371686 182898 371728 183134
rect 371408 182866 371728 182898
rect 371408 147454 371728 147486
rect 371408 147218 371450 147454
rect 371686 147218 371728 147454
rect 371408 147134 371728 147218
rect 371408 146898 371450 147134
rect 371686 146898 371728 147134
rect 371408 146866 371728 146898
rect 371408 111454 371728 111486
rect 371408 111218 371450 111454
rect 371686 111218 371728 111454
rect 371408 111134 371728 111218
rect 371408 110898 371450 111134
rect 371686 110898 371728 111134
rect 371408 110866 371728 110898
rect 371408 75454 371728 75486
rect 371408 75218 371450 75454
rect 371686 75218 371728 75454
rect 371408 75134 371728 75218
rect 371408 74898 371450 75134
rect 371686 74898 371728 75134
rect 371408 74866 371728 74898
rect 369234 46894 369854 58000
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 367691 40628 367757 40629
rect 367691 40564 367692 40628
rect 367756 40564 367757 40628
rect 367691 40563 367757 40564
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 58000
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 377262 2957 377322 539547
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 377259 2956 377325 2957
rect 377259 2892 377260 2956
rect 377324 2892 377325 2956
rect 377259 2891 377325 2892
rect 379794 -1306 380414 20898
rect 382230 8941 382290 539547
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 382227 8940 382293 8941
rect 382227 8876 382228 8940
rect 382292 8876 382293 8940
rect 382227 8875 382293 8876
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 -3226 384134 24618
rect 384990 18733 385050 539547
rect 386768 525454 387088 525486
rect 386768 525218 386810 525454
rect 387046 525218 387088 525454
rect 386768 525134 387088 525218
rect 386768 524898 386810 525134
rect 387046 524898 387088 525134
rect 386768 524866 387088 524898
rect 386768 489454 387088 489486
rect 386768 489218 386810 489454
rect 387046 489218 387088 489454
rect 386768 489134 387088 489218
rect 386768 488898 386810 489134
rect 387046 488898 387088 489134
rect 386768 488866 387088 488898
rect 386768 453454 387088 453486
rect 386768 453218 386810 453454
rect 387046 453218 387088 453454
rect 386768 453134 387088 453218
rect 386768 452898 386810 453134
rect 387046 452898 387088 453134
rect 386768 452866 387088 452898
rect 386768 417454 387088 417486
rect 386768 417218 386810 417454
rect 387046 417218 387088 417454
rect 386768 417134 387088 417218
rect 386768 416898 386810 417134
rect 387046 416898 387088 417134
rect 386768 416866 387088 416898
rect 386768 381454 387088 381486
rect 386768 381218 386810 381454
rect 387046 381218 387088 381454
rect 386768 381134 387088 381218
rect 386768 380898 386810 381134
rect 387046 380898 387088 381134
rect 386768 380866 387088 380898
rect 386768 345454 387088 345486
rect 386768 345218 386810 345454
rect 387046 345218 387088 345454
rect 386768 345134 387088 345218
rect 386768 344898 386810 345134
rect 387046 344898 387088 345134
rect 386768 344866 387088 344898
rect 386768 309454 387088 309486
rect 386768 309218 386810 309454
rect 387046 309218 387088 309454
rect 386768 309134 387088 309218
rect 386768 308898 386810 309134
rect 387046 308898 387088 309134
rect 386768 308866 387088 308898
rect 386768 273454 387088 273486
rect 386768 273218 386810 273454
rect 387046 273218 387088 273454
rect 386768 273134 387088 273218
rect 386768 272898 386810 273134
rect 387046 272898 387088 273134
rect 386768 272866 387088 272898
rect 386768 237454 387088 237486
rect 386768 237218 386810 237454
rect 387046 237218 387088 237454
rect 386768 237134 387088 237218
rect 386768 236898 386810 237134
rect 387046 236898 387088 237134
rect 386768 236866 387088 236898
rect 386768 201454 387088 201486
rect 386768 201218 386810 201454
rect 387046 201218 387088 201454
rect 386768 201134 387088 201218
rect 386768 200898 386810 201134
rect 387046 200898 387088 201134
rect 386768 200866 387088 200898
rect 386768 165454 387088 165486
rect 386768 165218 386810 165454
rect 387046 165218 387088 165454
rect 386768 165134 387088 165218
rect 386768 164898 386810 165134
rect 387046 164898 387088 165134
rect 386768 164866 387088 164898
rect 386768 129454 387088 129486
rect 386768 129218 386810 129454
rect 387046 129218 387088 129454
rect 386768 129134 387088 129218
rect 386768 128898 386810 129134
rect 387046 128898 387088 129134
rect 386768 128866 387088 128898
rect 386768 93454 387088 93486
rect 386768 93218 386810 93454
rect 387046 93218 387088 93454
rect 386768 93134 387088 93218
rect 386768 92898 386810 93134
rect 387046 92898 387088 93134
rect 386768 92866 387088 92898
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 384987 18732 385053 18733
rect 384987 18668 384988 18732
rect 385052 18668 385053 18732
rect 384987 18667 385053 18668
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 28338
rect 387934 24170 387994 539547
rect 388115 24172 388181 24173
rect 388115 24170 388116 24172
rect 387934 24110 388116 24170
rect 388115 24108 388116 24110
rect 388180 24108 388181 24172
rect 388115 24107 388181 24108
rect 389774 9077 389834 542539
rect 390954 542000 391574 572058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 542000 398414 542898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 542000 402134 546618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 542000 405854 550338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 542000 409574 554058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 542000 416414 560898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 542000 420134 564618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 542000 423854 568338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 542000 427574 572058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 542000 434414 542898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 542000 438134 546618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 542000 441854 550338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 393819 539612 393885 539613
rect 393819 539548 393820 539612
rect 393884 539548 393885 539612
rect 393819 539547 393885 539548
rect 400811 539612 400877 539613
rect 400811 539548 400812 539612
rect 400876 539548 400877 539612
rect 400811 539547 400877 539548
rect 393454 301018 393514 303502
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 389771 9076 389837 9077
rect 389771 9012 389772 9076
rect 389836 9012 389837 9076
rect 389771 9011 389837 9012
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 393822 4045 393882 539547
rect 397794 39454 398414 58000
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 393819 4044 393885 4045
rect 393819 3980 393820 4044
rect 393884 3980 393885 4044
rect 393819 3979 393885 3980
rect 397794 3454 398414 38898
rect 400814 13021 400874 539547
rect 417488 525454 417808 525486
rect 417488 525218 417530 525454
rect 417766 525218 417808 525454
rect 417488 525134 417808 525218
rect 417488 524898 417530 525134
rect 417766 524898 417808 525134
rect 417488 524866 417808 524898
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 402128 507454 402448 507486
rect 402128 507218 402170 507454
rect 402406 507218 402448 507454
rect 402128 507134 402448 507218
rect 402128 506898 402170 507134
rect 402406 506898 402448 507134
rect 402128 506866 402448 506898
rect 432848 507454 433168 507486
rect 432848 507218 432890 507454
rect 433126 507218 433168 507454
rect 432848 507134 433168 507218
rect 432848 506898 432890 507134
rect 433126 506898 433168 507134
rect 432848 506866 433168 506898
rect 417488 489454 417808 489486
rect 417488 489218 417530 489454
rect 417766 489218 417808 489454
rect 417488 489134 417808 489218
rect 417488 488898 417530 489134
rect 417766 488898 417808 489134
rect 417488 488866 417808 488898
rect 439451 488612 439517 488613
rect 439451 488548 439452 488612
rect 439516 488548 439517 488612
rect 439451 488547 439517 488548
rect 439454 488018 439514 488547
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 402128 471454 402448 471486
rect 402128 471218 402170 471454
rect 402406 471218 402448 471454
rect 402128 471134 402448 471218
rect 402128 470898 402170 471134
rect 402406 470898 402448 471134
rect 402128 470866 402448 470898
rect 432848 471454 433168 471486
rect 432848 471218 432890 471454
rect 433126 471218 433168 471454
rect 432848 471134 433168 471218
rect 432848 470898 432890 471134
rect 433126 470898 433168 471134
rect 432848 470866 433168 470898
rect 417488 453454 417808 453486
rect 417488 453218 417530 453454
rect 417766 453218 417808 453454
rect 417488 453134 417808 453218
rect 417488 452898 417530 453134
rect 417766 452898 417808 453134
rect 417488 452866 417808 452898
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 402128 435454 402448 435486
rect 402128 435218 402170 435454
rect 402406 435218 402448 435454
rect 402128 435134 402448 435218
rect 402128 434898 402170 435134
rect 402406 434898 402448 435134
rect 402128 434866 402448 434898
rect 432848 435454 433168 435486
rect 432848 435218 432890 435454
rect 433126 435218 433168 435454
rect 432848 435134 433168 435218
rect 432848 434898 432890 435134
rect 433126 434898 433168 435134
rect 432848 434866 433168 434898
rect 439270 425781 439330 425902
rect 439267 425780 439333 425781
rect 439267 425716 439268 425780
rect 439332 425716 439333 425780
rect 439267 425715 439333 425716
rect 417488 417454 417808 417486
rect 417488 417218 417530 417454
rect 417766 417218 417808 417454
rect 417488 417134 417808 417218
rect 417488 416898 417530 417134
rect 417766 416898 417808 417134
rect 417488 416866 417808 416898
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 402128 399454 402448 399486
rect 402128 399218 402170 399454
rect 402406 399218 402448 399454
rect 402128 399134 402448 399218
rect 402128 398898 402170 399134
rect 402406 398898 402448 399134
rect 402128 398866 402448 398898
rect 432848 399454 433168 399486
rect 432848 399218 432890 399454
rect 433126 399218 433168 399454
rect 432848 399134 433168 399218
rect 432848 398898 432890 399134
rect 433126 398898 433168 399134
rect 432848 398866 433168 398898
rect 439451 398172 439517 398173
rect 439451 398108 439452 398172
rect 439516 398108 439517 398172
rect 439451 398107 439517 398108
rect 439454 397578 439514 398107
rect 439451 392732 439517 392733
rect 439451 392668 439452 392732
rect 439516 392668 439517 392732
rect 439451 392667 439517 392668
rect 439454 391458 439514 392667
rect 417488 381454 417808 381486
rect 417488 381218 417530 381454
rect 417766 381218 417808 381454
rect 417488 381134 417808 381218
rect 417488 380898 417530 381134
rect 417766 380898 417808 381134
rect 417488 380866 417808 380898
rect 444954 374614 445574 410058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 453254 418301 453314 485742
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 453251 418300 453317 418301
rect 453251 418236 453252 418300
rect 453316 418236 453317 418300
rect 453251 418235 453317 418236
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 450491 404428 450557 404429
rect 450491 404364 450492 404428
rect 450556 404364 450557 404428
rect 450491 404363 450557 404364
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 402128 363454 402448 363486
rect 402128 363218 402170 363454
rect 402406 363218 402448 363454
rect 402128 363134 402448 363218
rect 402128 362898 402170 363134
rect 402406 362898 402448 363134
rect 402128 362866 402448 362898
rect 432848 363454 433168 363486
rect 432848 363218 432890 363454
rect 433126 363218 433168 363454
rect 432848 363134 433168 363218
rect 432848 362898 432890 363134
rect 433126 362898 433168 363134
rect 432848 362866 433168 362898
rect 439451 347308 439517 347309
rect 439451 347258 439452 347308
rect 439516 347258 439517 347308
rect 417488 345454 417808 345486
rect 417488 345218 417530 345454
rect 417766 345218 417808 345454
rect 417488 345134 417808 345218
rect 417488 344898 417530 345134
rect 417766 344898 417808 345134
rect 417488 344866 417808 344898
rect 444954 338614 445574 374058
rect 450494 343858 450554 404363
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 402128 327454 402448 327486
rect 402128 327218 402170 327454
rect 402406 327218 402448 327454
rect 402128 327134 402448 327218
rect 402128 326898 402170 327134
rect 402406 326898 402448 327134
rect 402128 326866 402448 326898
rect 432848 327454 433168 327486
rect 432848 327218 432890 327454
rect 433126 327218 433168 327454
rect 432848 327134 433168 327218
rect 432848 326898 432890 327134
rect 433126 326898 433168 327134
rect 432848 326866 433168 326898
rect 417488 309454 417808 309486
rect 417488 309218 417530 309454
rect 417766 309218 417808 309454
rect 417488 309134 417808 309218
rect 417488 308898 417530 309134
rect 417766 308898 417808 309134
rect 417488 308866 417808 308898
rect 422526 301018 422586 303502
rect 439454 302157 439514 303502
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 439451 302156 439517 302157
rect 439451 302092 439452 302156
rect 439516 302092 439517 302156
rect 439451 302091 439517 302092
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 449939 302156 450005 302157
rect 449939 302092 449940 302156
rect 450004 302092 450005 302156
rect 449939 302091 450005 302092
rect 402128 291454 402448 291486
rect 402128 291218 402170 291454
rect 402406 291218 402448 291454
rect 402128 291134 402448 291218
rect 402128 290898 402170 291134
rect 402406 290898 402448 291134
rect 402128 290866 402448 290898
rect 432848 291454 433168 291486
rect 432848 291218 432890 291454
rect 433126 291218 433168 291454
rect 432848 291134 433168 291218
rect 432848 290898 432890 291134
rect 433126 290898 433168 291134
rect 432848 290866 433168 290898
rect 417488 273454 417808 273486
rect 417488 273218 417530 273454
rect 417766 273218 417808 273454
rect 417488 273134 417808 273218
rect 417488 272898 417530 273134
rect 417766 272898 417808 273134
rect 417488 272866 417808 272898
rect 444954 266614 445574 302058
rect 449942 298213 450002 302091
rect 449939 298212 450005 298213
rect 449939 298148 449940 298212
rect 450004 298148 450005 298212
rect 449939 298147 450005 298148
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 402128 255454 402448 255486
rect 402128 255218 402170 255454
rect 402406 255218 402448 255454
rect 402128 255134 402448 255218
rect 402128 254898 402170 255134
rect 402406 254898 402448 255134
rect 402128 254866 402448 254898
rect 432848 255454 433168 255486
rect 432848 255218 432890 255454
rect 433126 255218 433168 255454
rect 432848 255134 433168 255218
rect 432848 254898 432890 255134
rect 433126 254898 433168 255134
rect 432848 254866 433168 254898
rect 417488 237454 417808 237486
rect 417488 237218 417530 237454
rect 417766 237218 417808 237454
rect 417488 237134 417808 237218
rect 417488 236898 417530 237134
rect 417766 236898 417808 237134
rect 417488 236866 417808 236898
rect 444954 230614 445574 266058
rect 451794 273454 452414 308898
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 450491 231980 450557 231981
rect 450491 231916 450492 231980
rect 450556 231916 450557 231980
rect 450491 231915 450557 231916
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 402128 219454 402448 219486
rect 402128 219218 402170 219454
rect 402406 219218 402448 219454
rect 402128 219134 402448 219218
rect 402128 218898 402170 219134
rect 402406 218898 402448 219134
rect 402128 218866 402448 218898
rect 432848 219454 433168 219486
rect 432848 219218 432890 219454
rect 433126 219218 433168 219454
rect 432848 219134 433168 219218
rect 432848 218898 432890 219134
rect 433126 218898 433168 219134
rect 432848 218866 433168 218898
rect 417488 201454 417808 201486
rect 417488 201218 417530 201454
rect 417766 201218 417808 201454
rect 417488 201134 417808 201218
rect 417488 200898 417530 201134
rect 417766 200898 417808 201134
rect 417488 200866 417808 200898
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 402128 183454 402448 183486
rect 402128 183218 402170 183454
rect 402406 183218 402448 183454
rect 402128 183134 402448 183218
rect 402128 182898 402170 183134
rect 402406 182898 402448 183134
rect 402128 182866 402448 182898
rect 432848 183454 433168 183486
rect 432848 183218 432890 183454
rect 433126 183218 433168 183454
rect 432848 183134 433168 183218
rect 432848 182898 432890 183134
rect 433126 182898 433168 183134
rect 432848 182866 433168 182898
rect 417488 165454 417808 165486
rect 417488 165218 417530 165454
rect 417766 165218 417808 165454
rect 417488 165134 417808 165218
rect 417488 164898 417530 165134
rect 417766 164898 417808 165134
rect 417488 164866 417808 164898
rect 444954 158614 445574 194058
rect 450494 179298 450554 231915
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 402128 147454 402448 147486
rect 402128 147218 402170 147454
rect 402406 147218 402448 147454
rect 402128 147134 402448 147218
rect 402128 146898 402170 147134
rect 402406 146898 402448 147134
rect 402128 146866 402448 146898
rect 432848 147454 433168 147486
rect 432848 147218 432890 147454
rect 433126 147218 433168 147454
rect 432848 147134 433168 147218
rect 432848 146898 432890 147134
rect 433126 146898 433168 147134
rect 432848 146866 433168 146898
rect 417488 129454 417808 129486
rect 417488 129218 417530 129454
rect 417766 129218 417808 129454
rect 417488 129134 417808 129218
rect 417488 128898 417530 129134
rect 417766 128898 417808 129134
rect 417488 128866 417808 128898
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 402128 111454 402448 111486
rect 402128 111218 402170 111454
rect 402406 111218 402448 111454
rect 402128 111134 402448 111218
rect 402128 110898 402170 111134
rect 402406 110898 402448 111134
rect 402128 110866 402448 110898
rect 432848 111454 433168 111486
rect 432848 111218 432890 111454
rect 433126 111218 433168 111454
rect 432848 111134 433168 111218
rect 432848 110898 432890 111134
rect 433126 110898 433168 111134
rect 432848 110866 433168 110898
rect 417488 93454 417808 93486
rect 417488 93218 417530 93454
rect 417766 93218 417808 93454
rect 417488 93134 417808 93218
rect 417488 92898 417530 93134
rect 417766 92898 417808 93134
rect 417488 92866 417808 92898
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 402128 75454 402448 75486
rect 402128 75218 402170 75454
rect 402406 75218 402448 75454
rect 402128 75134 402448 75218
rect 402128 74898 402170 75134
rect 402406 74898 402448 75134
rect 402128 74866 402448 74898
rect 432848 75454 433168 75486
rect 432848 75218 432890 75454
rect 433126 75218 433168 75454
rect 432848 75134 433168 75218
rect 432848 74898 432890 75134
rect 433126 74898 433168 75134
rect 432848 74866 433168 74898
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 400811 13020 400877 13021
rect 400811 12956 400812 13020
rect 400876 12956 400877 13020
rect 400811 12955 400877 12956
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 453254 138141 453314 274262
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 453251 138140 453317 138141
rect 453251 138076 453252 138140
rect 453316 138076 453317 138140
rect 453251 138075 453317 138076
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 471099 311948 471165 311949
rect 471099 311884 471100 311948
rect 471164 311884 471165 311948
rect 471099 311883 471165 311884
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 468342 125629 468402 213062
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 471102 160938 471162 311883
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 468339 125628 468405 125629
rect 468339 125564 468340 125628
rect 468404 125564 468405 125628
rect 468339 125563 468405 125564
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 500171 378180 500237 378181
rect 500171 378116 500172 378180
rect 500236 378116 500237 378180
rect 500171 378115 500237 378116
rect 500174 371738 500234 378115
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 21134 425902 21370 426138
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 22606 397342 22842 397578
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 34934 487782 35170 488018
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 32174 391222 32410 391458
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 33646 347022 33882 347258
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 36406 433382 36642 433618
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 60510 485892 60746 485978
rect 60510 485828 60596 485892
rect 60596 485828 60660 485892
rect 60660 485828 60746 485892
rect 60510 485742 60746 485828
rect 64250 471218 64486 471454
rect 64250 470898 64486 471134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 64250 435218 64486 435454
rect 64250 434898 64486 435134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 64250 399218 64486 399454
rect 64250 398898 64486 399134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 60510 371502 60746 371738
rect 64250 363218 64486 363454
rect 64250 362898 64486 363134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 60510 343772 60746 343858
rect 60510 343708 60596 343772
rect 60596 343708 60660 343772
rect 60660 343708 60746 343772
rect 60510 343622 60746 343708
rect 64250 327218 64486 327454
rect 64250 326898 64486 327134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 60510 303502 60746 303738
rect 65294 303502 65530 303738
rect 65294 300782 65530 301018
rect 64250 291218 64486 291454
rect 64250 290898 64486 291134
rect 60510 274484 60596 274498
rect 60596 274484 60660 274498
rect 60660 274484 60746 274498
rect 60510 274262 60746 274484
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 64250 255218 64486 255454
rect 64250 254898 64486 255134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 64250 219218 64486 219454
rect 64250 218898 64486 219134
rect 60510 213212 60746 213298
rect 60510 213148 60596 213212
rect 60596 213148 60660 213212
rect 60660 213148 60746 213212
rect 60510 213062 60746 213148
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 64250 183218 64486 183454
rect 64250 182898 64486 183134
rect 60510 179284 60596 179298
rect 60596 179284 60660 179298
rect 60660 179284 60746 179298
rect 60510 179062 60746 179284
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 60510 160852 60746 160938
rect 60510 160788 60596 160852
rect 60596 160788 60660 160852
rect 60660 160788 60746 160852
rect 60510 160702 60746 160788
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 64250 111218 64486 111454
rect 64250 110898 64486 111134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 64250 75218 64486 75454
rect 64250 74898 64486 75134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 61982 4302 62218 4538
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 79610 525218 79846 525454
rect 79610 524898 79846 525134
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 79610 489218 79846 489454
rect 79610 488898 79846 489134
rect 94970 471218 95206 471454
rect 94970 470898 95206 471134
rect 79610 453218 79846 453454
rect 79610 452898 79846 453134
rect 94970 435218 95206 435454
rect 94970 434898 95206 435134
rect 79610 417218 79846 417454
rect 79610 416898 79846 417134
rect 94970 399218 95206 399454
rect 94970 398898 95206 399134
rect 79610 381218 79846 381454
rect 79610 380898 79846 381134
rect 94970 363218 95206 363454
rect 94970 362898 95206 363134
rect 79610 345218 79846 345454
rect 79610 344898 79846 345134
rect 94970 327218 95206 327454
rect 94970 326898 95206 327134
rect 79610 309218 79846 309454
rect 79610 308898 79846 309134
rect 85350 303502 85586 303738
rect 93814 303502 94050 303738
rect 85350 300782 85586 301018
rect 93814 300782 94050 301018
rect 94970 291218 95206 291454
rect 94970 290898 95206 291134
rect 79610 273218 79846 273454
rect 79610 272898 79846 273134
rect 94970 255218 95206 255454
rect 94970 254898 95206 255134
rect 79610 237218 79846 237454
rect 79610 236898 79846 237134
rect 94970 219218 95206 219454
rect 94970 218898 95206 219134
rect 79610 201218 79846 201454
rect 79610 200898 79846 201134
rect 94970 183218 95206 183454
rect 94970 182898 95206 183134
rect 79610 165218 79846 165454
rect 79610 164898 79846 165134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 79610 129218 79846 129454
rect 79610 128898 79846 129134
rect 94970 111218 95206 111454
rect 94970 110898 95206 111134
rect 79610 93218 79846 93454
rect 79610 92898 79846 93134
rect 94970 75218 95206 75454
rect 94970 74898 95206 75134
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 110330 525218 110566 525454
rect 110330 524898 110566 525134
rect 110330 489218 110566 489454
rect 110330 488898 110566 489134
rect 110330 453218 110566 453454
rect 110330 452898 110566 453134
rect 110330 417218 110566 417454
rect 110330 416898 110566 417134
rect 110330 381218 110566 381454
rect 110330 380898 110566 381134
rect 110330 345218 110566 345454
rect 110330 344898 110566 345134
rect 110330 309218 110566 309454
rect 110330 308898 110566 309134
rect 113686 303502 113922 303738
rect 113686 300782 113922 301018
rect 110330 273218 110566 273454
rect 110330 272898 110566 273134
rect 110330 237218 110566 237454
rect 110330 236898 110566 237134
rect 110330 201218 110566 201454
rect 110330 200898 110566 201134
rect 110330 165218 110566 165454
rect 110330 164898 110566 165134
rect 110330 129218 110566 129454
rect 110330 128898 110566 129134
rect 110330 93218 110566 93454
rect 110330 92898 110566 93134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 125690 471218 125926 471454
rect 125690 470898 125926 471134
rect 125690 435218 125926 435454
rect 125690 434898 125926 435134
rect 125690 399218 125926 399454
rect 125690 398898 125926 399134
rect 125690 363218 125926 363454
rect 125690 362898 125926 363134
rect 125690 327218 125926 327454
rect 125690 326898 125926 327134
rect 125690 291218 125926 291454
rect 125690 290898 125926 291134
rect 125690 255218 125926 255454
rect 125690 254898 125926 255134
rect 125690 219218 125926 219454
rect 125690 218898 125926 219134
rect 125690 183218 125926 183454
rect 125690 182898 125926 183134
rect 125690 147218 125926 147454
rect 125690 146898 125926 147134
rect 125690 111218 125926 111454
rect 125690 110898 125926 111134
rect 125690 75218 125926 75454
rect 125690 74898 125926 75134
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 141050 525218 141286 525454
rect 141050 524898 141286 525134
rect 141050 489218 141286 489454
rect 141050 488898 141286 489134
rect 141050 453218 141286 453454
rect 141050 452898 141286 453134
rect 141050 417218 141286 417454
rect 141050 416898 141286 417134
rect 141050 381218 141286 381454
rect 141050 380898 141286 381134
rect 141050 345218 141286 345454
rect 141050 344898 141286 345134
rect 141050 309218 141286 309454
rect 141050 308898 141286 309134
rect 142942 303502 143178 303738
rect 142942 300782 143178 301018
rect 141050 273218 141286 273454
rect 141050 272898 141286 273134
rect 141050 237218 141286 237454
rect 141050 236898 141286 237134
rect 141050 201218 141286 201454
rect 141050 200898 141286 201134
rect 141050 165218 141286 165454
rect 141050 164898 141286 165134
rect 141050 129218 141286 129454
rect 141050 128898 141286 129134
rect 141050 93218 141286 93454
rect 141050 92898 141286 93134
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 153798 303502 154034 303738
rect 153798 300782 154034 301018
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 156410 471218 156646 471454
rect 156410 470898 156646 471134
rect 156410 435218 156646 435454
rect 156410 434898 156646 435134
rect 156410 399218 156646 399454
rect 156410 398898 156646 399134
rect 156410 363218 156646 363454
rect 156410 362898 156646 363134
rect 156410 327218 156646 327454
rect 156410 326898 156646 327134
rect 161526 303502 161762 303738
rect 161526 300782 161762 301018
rect 156410 291218 156646 291454
rect 156410 290898 156646 291134
rect 156410 255218 156646 255454
rect 156410 254898 156646 255134
rect 156410 219218 156646 219454
rect 156410 218898 156646 219134
rect 156410 183218 156646 183454
rect 156410 182898 156646 183134
rect 156410 147218 156646 147454
rect 156410 146898 156646 147134
rect 156410 111218 156646 111454
rect 156410 110898 156646 111134
rect 156410 75218 156646 75454
rect 156410 74898 156646 75134
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 171770 525218 172006 525454
rect 171770 524898 172006 525134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 171770 489218 172006 489454
rect 171770 488898 172006 489134
rect 187130 471218 187366 471454
rect 187130 470898 187366 471134
rect 171770 453218 172006 453454
rect 171770 452898 172006 453134
rect 187130 435218 187366 435454
rect 187130 434898 187366 435134
rect 171770 417218 172006 417454
rect 171770 416898 172006 417134
rect 187130 399218 187366 399454
rect 187130 398898 187366 399134
rect 171770 381218 172006 381454
rect 171770 380898 172006 381134
rect 187130 363218 187366 363454
rect 187130 362898 187366 363134
rect 171770 345218 172006 345454
rect 171770 344898 172006 345134
rect 187130 327218 187366 327454
rect 187130 326898 187366 327134
rect 171770 309218 172006 309454
rect 171770 308898 172006 309134
rect 190598 303502 190834 303738
rect 190598 300782 190834 301018
rect 187130 291218 187366 291454
rect 187130 290898 187366 291134
rect 171770 273218 172006 273454
rect 171770 272898 172006 273134
rect 187130 255218 187366 255454
rect 187130 254898 187366 255134
rect 171770 237218 172006 237454
rect 171770 236898 172006 237134
rect 187130 219218 187366 219454
rect 187130 218898 187366 219134
rect 171770 201218 172006 201454
rect 171770 200898 172006 201134
rect 187130 183218 187366 183454
rect 187130 182898 187366 183134
rect 171770 165218 172006 165454
rect 171770 164898 172006 165134
rect 187130 147218 187366 147454
rect 187130 146898 187366 147134
rect 171770 129218 172006 129454
rect 171770 128898 172006 129134
rect 187130 111218 187366 111454
rect 187130 110898 187366 111134
rect 171770 93218 172006 93454
rect 171770 92898 172006 93134
rect 187130 75218 187366 75454
rect 187130 74898 187366 75134
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 202490 525218 202726 525454
rect 202490 524898 202726 525134
rect 202490 489218 202726 489454
rect 202490 488898 202726 489134
rect 202490 453218 202726 453454
rect 202490 452898 202726 453134
rect 202490 417218 202726 417454
rect 202490 416898 202726 417134
rect 202490 381218 202726 381454
rect 202490 380898 202726 381134
rect 202490 345218 202726 345454
rect 202490 344898 202726 345134
rect 202490 309218 202726 309454
rect 202490 308898 202726 309134
rect 202490 273218 202726 273454
rect 202490 272898 202726 273134
rect 202490 237218 202726 237454
rect 202490 236898 202726 237134
rect 202490 201218 202726 201454
rect 202490 200898 202726 201134
rect 202490 165218 202726 165454
rect 202490 164898 202726 165134
rect 202490 129218 202726 129454
rect 202490 128898 202726 129134
rect 202490 93218 202726 93454
rect 202490 92898 202726 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 217850 471218 218086 471454
rect 217850 470898 218086 471134
rect 217850 435218 218086 435454
rect 217850 434898 218086 435134
rect 217850 399218 218086 399454
rect 217850 398898 218086 399134
rect 217850 363218 218086 363454
rect 217850 362898 218086 363134
rect 217850 327218 218086 327454
rect 217850 326898 218086 327134
rect 211206 303502 211442 303738
rect 211206 300782 211442 301018
rect 217850 291218 218086 291454
rect 217850 290898 218086 291134
rect 217850 255218 218086 255454
rect 217850 254898 218086 255134
rect 217850 219218 218086 219454
rect 217850 218898 218086 219134
rect 217850 183218 218086 183454
rect 217850 182898 218086 183134
rect 217850 147218 218086 147454
rect 217850 146898 218086 147134
rect 217850 111218 218086 111454
rect 217850 110898 218086 111134
rect 217850 75218 218086 75454
rect 217850 74898 218086 75134
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 220222 303502 220458 303738
rect 220222 300782 220458 301018
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 233210 525218 233446 525454
rect 233210 524898 233446 525134
rect 233210 489218 233446 489454
rect 233210 488898 233446 489134
rect 233210 453218 233446 453454
rect 233210 452898 233446 453134
rect 233210 417218 233446 417454
rect 233210 416898 233446 417134
rect 233210 381218 233446 381454
rect 233210 380898 233446 381134
rect 233210 345218 233446 345454
rect 233210 344898 233446 345134
rect 233210 309218 233446 309454
rect 233210 308898 233446 309134
rect 233210 273218 233446 273454
rect 233210 272898 233446 273134
rect 233210 237218 233446 237454
rect 233210 236898 233446 237134
rect 233210 201218 233446 201454
rect 233210 200898 233446 201134
rect 233210 165218 233446 165454
rect 233210 164898 233446 165134
rect 233210 129218 233446 129454
rect 233210 128898 233446 129134
rect 233210 93218 233446 93454
rect 233210 92898 233446 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 248570 471218 248806 471454
rect 248570 470898 248806 471134
rect 248570 435218 248806 435454
rect 248570 434898 248806 435134
rect 248570 399218 248806 399454
rect 248570 398898 248806 399134
rect 248570 363218 248806 363454
rect 248570 362898 248806 363134
rect 248570 327218 248806 327454
rect 248570 326898 248806 327134
rect 249294 303502 249530 303738
rect 249294 300782 249530 301018
rect 248570 291218 248806 291454
rect 248570 290898 248806 291134
rect 248570 255218 248806 255454
rect 248570 254898 248806 255134
rect 248570 219218 248806 219454
rect 248570 218898 248806 219134
rect 248570 183218 248806 183454
rect 248570 182898 248806 183134
rect 248570 147218 248806 147454
rect 248570 146898 248806 147134
rect 248570 111218 248806 111454
rect 248570 110898 248806 111134
rect 248570 75218 248806 75454
rect 248570 74898 248806 75134
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 263930 525218 264166 525454
rect 263930 524898 264166 525134
rect 263930 489218 264166 489454
rect 263930 488898 264166 489134
rect 263930 453218 264166 453454
rect 263930 452898 264166 453134
rect 263930 417218 264166 417454
rect 263930 416898 264166 417134
rect 263930 381218 264166 381454
rect 263930 380898 264166 381134
rect 263930 345218 264166 345454
rect 263930 344898 264166 345134
rect 263930 309218 264166 309454
rect 263930 308898 264166 309134
rect 263930 273218 264166 273454
rect 263930 272898 264166 273134
rect 263930 237218 264166 237454
rect 263930 236898 264166 237134
rect 263930 201218 264166 201454
rect 263930 200898 264166 201134
rect 263930 165218 264166 165454
rect 263930 164898 264166 165134
rect 263930 129218 264166 129454
rect 263930 128898 264166 129134
rect 263930 93218 264166 93454
rect 263930 92898 264166 93134
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 267878 303502 268114 303738
rect 267878 300782 268114 301018
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 279290 471218 279526 471454
rect 279290 470898 279526 471134
rect 279290 435218 279526 435454
rect 279290 434898 279526 435134
rect 279290 399218 279526 399454
rect 279290 398898 279526 399134
rect 279290 363218 279526 363454
rect 279290 362898 279526 363134
rect 279290 327218 279526 327454
rect 279290 326898 279526 327134
rect 279290 291218 279526 291454
rect 279290 290898 279526 291134
rect 279290 255218 279526 255454
rect 279290 254898 279526 255134
rect 279290 219218 279526 219454
rect 279290 218898 279526 219134
rect 279290 183218 279526 183454
rect 279290 182898 279526 183134
rect 279290 147218 279526 147454
rect 279290 146898 279526 147134
rect 279290 111218 279526 111454
rect 279290 110898 279526 111134
rect 279290 75218 279526 75454
rect 279290 74898 279526 75134
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 294650 525218 294886 525454
rect 294650 524898 294886 525134
rect 294650 489218 294886 489454
rect 294650 488898 294886 489134
rect 294650 453218 294886 453454
rect 294650 452898 294886 453134
rect 294650 417218 294886 417454
rect 294650 416898 294886 417134
rect 294650 381218 294886 381454
rect 294650 380898 294886 381134
rect 294650 345218 294886 345454
rect 294650 344898 294886 345134
rect 294650 309218 294886 309454
rect 294650 308898 294886 309134
rect 287566 303502 287802 303738
rect 287566 300782 287802 301018
rect 294650 273218 294886 273454
rect 294650 272898 294886 273134
rect 294650 237218 294886 237454
rect 294650 236898 294886 237134
rect 294650 201218 294886 201454
rect 294650 200898 294886 201134
rect 294650 165218 294886 165454
rect 294650 164898 294886 165134
rect 294650 129218 294886 129454
rect 294650 128898 294886 129134
rect 294650 93218 294886 93454
rect 294650 92898 294886 93134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 310010 507218 310246 507454
rect 310010 506898 310246 507134
rect 310010 471218 310246 471454
rect 310010 470898 310246 471134
rect 310010 435218 310246 435454
rect 310010 434898 310246 435134
rect 310010 399218 310246 399454
rect 310010 398898 310246 399134
rect 310010 363218 310246 363454
rect 310010 362898 310246 363134
rect 310010 327218 310246 327454
rect 310010 326898 310246 327134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 310010 291218 310246 291454
rect 310010 290898 310246 291134
rect 310010 255218 310246 255454
rect 310010 254898 310246 255134
rect 310010 219218 310246 219454
rect 310010 218898 310246 219134
rect 310010 183218 310246 183454
rect 310010 182898 310246 183134
rect 310010 147218 310246 147454
rect 310010 146898 310246 147134
rect 310010 111218 310246 111454
rect 310010 110898 310246 111134
rect 310010 75218 310246 75454
rect 310010 74898 310246 75134
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 309094 4302 309330 4538
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 316454 303502 316690 303738
rect 316454 300782 316690 301018
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325370 525218 325606 525454
rect 325370 524898 325606 525134
rect 325370 489218 325606 489454
rect 325370 488898 325606 489134
rect 325370 453218 325606 453454
rect 325370 452898 325606 453134
rect 325370 417218 325606 417454
rect 325370 416898 325606 417134
rect 325370 381218 325606 381454
rect 325370 380898 325606 381134
rect 325370 345218 325606 345454
rect 325370 344898 325606 345134
rect 325370 309218 325606 309454
rect 325370 308898 325606 309134
rect 325370 273218 325606 273454
rect 325370 272898 325606 273134
rect 325370 237218 325606 237454
rect 325370 236898 325606 237134
rect 325370 201218 325606 201454
rect 325370 200898 325606 201134
rect 325370 165218 325606 165454
rect 325370 164898 325606 165134
rect 325370 129218 325606 129454
rect 325370 128898 325606 129134
rect 325370 93218 325606 93454
rect 325370 92898 325606 93134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 340730 507218 340966 507454
rect 340730 506898 340966 507134
rect 340730 471218 340966 471454
rect 340730 470898 340966 471134
rect 340730 435218 340966 435454
rect 340730 434898 340966 435134
rect 340730 399218 340966 399454
rect 340730 398898 340966 399134
rect 340730 363218 340966 363454
rect 340730 362898 340966 363134
rect 340730 327218 340966 327454
rect 340730 326898 340966 327134
rect 340730 291218 340966 291454
rect 340730 290898 340966 291134
rect 340730 255218 340966 255454
rect 340730 254898 340966 255134
rect 340730 219218 340966 219454
rect 340730 218898 340966 219134
rect 340730 183218 340966 183454
rect 340730 182898 340966 183134
rect 340730 147218 340966 147454
rect 340730 146898 340966 147134
rect 340730 111218 340966 111454
rect 340730 110898 340966 111134
rect 340730 75218 340966 75454
rect 340730 74898 340966 75134
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 356090 525218 356326 525454
rect 356090 524898 356326 525134
rect 356090 489218 356326 489454
rect 356090 488898 356326 489134
rect 356090 453218 356326 453454
rect 356090 452898 356326 453134
rect 356090 417218 356326 417454
rect 356090 416898 356326 417134
rect 356090 381218 356326 381454
rect 356090 380898 356326 381134
rect 356090 345218 356326 345454
rect 356090 344898 356326 345134
rect 356090 309218 356326 309454
rect 356090 308898 356326 309134
rect 354910 303502 355146 303738
rect 354910 300782 355146 301018
rect 356090 273218 356326 273454
rect 356090 272898 356326 273134
rect 356090 237218 356326 237454
rect 356090 236898 356326 237134
rect 356090 201218 356326 201454
rect 356090 200898 356326 201134
rect 356090 165218 356326 165454
rect 356090 164898 356326 165134
rect 356090 129218 356326 129454
rect 356090 128898 356326 129134
rect 356090 93218 356326 93454
rect 356090 92898 356326 93134
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 371450 507218 371686 507454
rect 371450 506898 371686 507134
rect 371450 471218 371686 471454
rect 371450 470898 371686 471134
rect 371450 435218 371686 435454
rect 371450 434898 371686 435134
rect 371450 399218 371686 399454
rect 371450 398898 371686 399134
rect 371450 363218 371686 363454
rect 371450 362898 371686 363134
rect 371450 327218 371686 327454
rect 371450 326898 371686 327134
rect 374046 303502 374282 303738
rect 374046 300782 374282 301018
rect 371450 291218 371686 291454
rect 371450 290898 371686 291134
rect 371450 255218 371686 255454
rect 371450 254898 371686 255134
rect 371450 219218 371686 219454
rect 371450 218898 371686 219134
rect 371450 183218 371686 183454
rect 371450 182898 371686 183134
rect 371450 147218 371686 147454
rect 371450 146898 371686 147134
rect 371450 111218 371686 111454
rect 371450 110898 371686 111134
rect 371450 75218 371686 75454
rect 371450 74898 371686 75134
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 386810 525218 387046 525454
rect 386810 524898 387046 525134
rect 386810 489218 387046 489454
rect 386810 488898 387046 489134
rect 386810 453218 387046 453454
rect 386810 452898 387046 453134
rect 386810 417218 387046 417454
rect 386810 416898 387046 417134
rect 386810 381218 387046 381454
rect 386810 380898 387046 381134
rect 386810 345218 387046 345454
rect 386810 344898 387046 345134
rect 386810 309218 387046 309454
rect 386810 308898 387046 309134
rect 386810 273218 387046 273454
rect 386810 272898 387046 273134
rect 386810 237218 387046 237454
rect 386810 236898 387046 237134
rect 386810 201218 387046 201454
rect 386810 200898 387046 201134
rect 386810 165218 387046 165454
rect 386810 164898 387046 165134
rect 386810 129218 387046 129454
rect 386810 128898 387046 129134
rect 386810 93218 387046 93454
rect 386810 92898 387046 93134
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 393366 303502 393602 303738
rect 393366 300782 393602 301018
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 417530 525218 417766 525454
rect 417530 524898 417766 525134
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 402170 507218 402406 507454
rect 402170 506898 402406 507134
rect 432890 507218 433126 507454
rect 432890 506898 433126 507134
rect 417530 489218 417766 489454
rect 417530 488898 417766 489134
rect 439366 487782 439602 488018
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 402170 471218 402406 471454
rect 402170 470898 402406 471134
rect 432890 471218 433126 471454
rect 432890 470898 433126 471134
rect 417530 453218 417766 453454
rect 417530 452898 417766 453134
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 402170 435218 402406 435454
rect 402170 434898 402406 435134
rect 432890 435218 433126 435454
rect 432890 434898 433126 435134
rect 439366 433532 439602 433618
rect 439366 433468 439452 433532
rect 439452 433468 439516 433532
rect 439516 433468 439602 433532
rect 439366 433382 439602 433468
rect 439182 425902 439418 426138
rect 417530 417218 417766 417454
rect 417530 416898 417766 417134
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 402170 399218 402406 399454
rect 402170 398898 402406 399134
rect 432890 399218 433126 399454
rect 432890 398898 433126 399134
rect 439366 397342 439602 397578
rect 439366 391222 439602 391458
rect 417530 381218 417766 381454
rect 417530 380898 417766 381134
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 453166 485742 453402 485978
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 402170 363218 402406 363454
rect 402170 362898 402406 363134
rect 432890 363218 433126 363454
rect 432890 362898 433126 363134
rect 439366 347244 439452 347258
rect 439452 347244 439516 347258
rect 439516 347244 439602 347258
rect 439366 347022 439602 347244
rect 417530 345218 417766 345454
rect 417530 344898 417766 345134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 450406 343622 450642 343858
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 402170 327218 402406 327454
rect 402170 326898 402406 327134
rect 432890 327218 433126 327454
rect 432890 326898 433126 327134
rect 417530 309218 417766 309454
rect 417530 308898 417766 309134
rect 422438 303502 422674 303738
rect 439366 303502 439602 303738
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 422438 300782 422674 301018
rect 402170 291218 402406 291454
rect 402170 290898 402406 291134
rect 432890 291218 433126 291454
rect 432890 290898 433126 291134
rect 417530 273218 417766 273454
rect 417530 272898 417766 273134
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 402170 255218 402406 255454
rect 402170 254898 402406 255134
rect 432890 255218 433126 255454
rect 432890 254898 433126 255134
rect 417530 237218 417766 237454
rect 417530 236898 417766 237134
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 453166 274262 453402 274498
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 402170 219218 402406 219454
rect 402170 218898 402406 219134
rect 432890 219218 433126 219454
rect 432890 218898 433126 219134
rect 417530 201218 417766 201454
rect 417530 200898 417766 201134
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 402170 183218 402406 183454
rect 402170 182898 402406 183134
rect 432890 183218 433126 183454
rect 432890 182898 433126 183134
rect 417530 165218 417766 165454
rect 417530 164898 417766 165134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 450406 179062 450642 179298
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 402170 147218 402406 147454
rect 402170 146898 402406 147134
rect 432890 147218 433126 147454
rect 432890 146898 433126 147134
rect 417530 129218 417766 129454
rect 417530 128898 417766 129134
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 402170 111218 402406 111454
rect 402170 110898 402406 111134
rect 432890 111218 433126 111454
rect 432890 110898 433126 111134
rect 417530 93218 417766 93454
rect 417530 92898 417766 93134
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 402170 75218 402406 75454
rect 402170 74898 402406 75134
rect 432890 75218 433126 75454
rect 432890 74898 433126 75134
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 468254 213062 468490 213298
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 471014 160702 471250 160938
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 500086 371502 500322 371738
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 79610 525454
rect 79846 525218 110330 525454
rect 110566 525218 141050 525454
rect 141286 525218 171770 525454
rect 172006 525218 202490 525454
rect 202726 525218 233210 525454
rect 233446 525218 263930 525454
rect 264166 525218 294650 525454
rect 294886 525218 325370 525454
rect 325606 525218 356090 525454
rect 356326 525218 386810 525454
rect 387046 525218 417530 525454
rect 417766 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 79610 525134
rect 79846 524898 110330 525134
rect 110566 524898 141050 525134
rect 141286 524898 171770 525134
rect 172006 524898 202490 525134
rect 202726 524898 233210 525134
rect 233446 524898 263930 525134
rect 264166 524898 294650 525134
rect 294886 524898 325370 525134
rect 325606 524898 356090 525134
rect 356326 524898 386810 525134
rect 387046 524898 417530 525134
rect 417766 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 310010 507454
rect 310246 507218 340730 507454
rect 340966 507218 371450 507454
rect 371686 507218 402170 507454
rect 402406 507218 432890 507454
rect 433126 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 310010 507134
rect 310246 506898 340730 507134
rect 340966 506898 371450 507134
rect 371686 506898 402170 507134
rect 402406 506898 432890 507134
rect 433126 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 79610 489454
rect 79846 489218 110330 489454
rect 110566 489218 141050 489454
rect 141286 489218 171770 489454
rect 172006 489218 202490 489454
rect 202726 489218 233210 489454
rect 233446 489218 263930 489454
rect 264166 489218 294650 489454
rect 294886 489218 325370 489454
rect 325606 489218 356090 489454
rect 356326 489218 386810 489454
rect 387046 489218 417530 489454
rect 417766 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 79610 489134
rect 79846 488898 110330 489134
rect 110566 488898 141050 489134
rect 141286 488898 171770 489134
rect 172006 488898 202490 489134
rect 202726 488898 233210 489134
rect 233446 488898 263930 489134
rect 264166 488898 294650 489134
rect 294886 488898 325370 489134
rect 325606 488898 356090 489134
rect 356326 488898 386810 489134
rect 387046 488898 417530 489134
rect 417766 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect 34892 488018 439644 488060
rect 34892 487782 34934 488018
rect 35170 487782 439366 488018
rect 439602 487782 439644 488018
rect 34892 487740 439644 487782
rect 60468 485978 453444 486020
rect 60468 485742 60510 485978
rect 60746 485742 453166 485978
rect 453402 485742 453444 485978
rect 60468 485700 453444 485742
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 64250 471454
rect 64486 471218 94970 471454
rect 95206 471218 125690 471454
rect 125926 471218 156410 471454
rect 156646 471218 187130 471454
rect 187366 471218 217850 471454
rect 218086 471218 248570 471454
rect 248806 471218 279290 471454
rect 279526 471218 310010 471454
rect 310246 471218 340730 471454
rect 340966 471218 371450 471454
rect 371686 471218 402170 471454
rect 402406 471218 432890 471454
rect 433126 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 64250 471134
rect 64486 470898 94970 471134
rect 95206 470898 125690 471134
rect 125926 470898 156410 471134
rect 156646 470898 187130 471134
rect 187366 470898 217850 471134
rect 218086 470898 248570 471134
rect 248806 470898 279290 471134
rect 279526 470898 310010 471134
rect 310246 470898 340730 471134
rect 340966 470898 371450 471134
rect 371686 470898 402170 471134
rect 402406 470898 432890 471134
rect 433126 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 79610 453454
rect 79846 453218 110330 453454
rect 110566 453218 141050 453454
rect 141286 453218 171770 453454
rect 172006 453218 202490 453454
rect 202726 453218 233210 453454
rect 233446 453218 263930 453454
rect 264166 453218 294650 453454
rect 294886 453218 325370 453454
rect 325606 453218 356090 453454
rect 356326 453218 386810 453454
rect 387046 453218 417530 453454
rect 417766 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 79610 453134
rect 79846 452898 110330 453134
rect 110566 452898 141050 453134
rect 141286 452898 171770 453134
rect 172006 452898 202490 453134
rect 202726 452898 233210 453134
rect 233446 452898 263930 453134
rect 264166 452898 294650 453134
rect 294886 452898 325370 453134
rect 325606 452898 356090 453134
rect 356326 452898 386810 453134
rect 387046 452898 417530 453134
rect 417766 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 64250 435454
rect 64486 435218 94970 435454
rect 95206 435218 125690 435454
rect 125926 435218 156410 435454
rect 156646 435218 187130 435454
rect 187366 435218 217850 435454
rect 218086 435218 248570 435454
rect 248806 435218 279290 435454
rect 279526 435218 310010 435454
rect 310246 435218 340730 435454
rect 340966 435218 371450 435454
rect 371686 435218 402170 435454
rect 402406 435218 432890 435454
rect 433126 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 64250 435134
rect 64486 434898 94970 435134
rect 95206 434898 125690 435134
rect 125926 434898 156410 435134
rect 156646 434898 187130 435134
rect 187366 434898 217850 435134
rect 218086 434898 248570 435134
rect 248806 434898 279290 435134
rect 279526 434898 310010 435134
rect 310246 434898 340730 435134
rect 340966 434898 371450 435134
rect 371686 434898 402170 435134
rect 402406 434898 432890 435134
rect 433126 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect 36364 433618 439644 433660
rect 36364 433382 36406 433618
rect 36642 433382 439366 433618
rect 439602 433382 439644 433618
rect 36364 433340 439644 433382
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect 21092 426138 439460 426180
rect 21092 425902 21134 426138
rect 21370 425902 439182 426138
rect 439418 425902 439460 426138
rect 21092 425860 439460 425902
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 79610 417454
rect 79846 417218 110330 417454
rect 110566 417218 141050 417454
rect 141286 417218 171770 417454
rect 172006 417218 202490 417454
rect 202726 417218 233210 417454
rect 233446 417218 263930 417454
rect 264166 417218 294650 417454
rect 294886 417218 325370 417454
rect 325606 417218 356090 417454
rect 356326 417218 386810 417454
rect 387046 417218 417530 417454
rect 417766 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 79610 417134
rect 79846 416898 110330 417134
rect 110566 416898 141050 417134
rect 141286 416898 171770 417134
rect 172006 416898 202490 417134
rect 202726 416898 233210 417134
rect 233446 416898 263930 417134
rect 264166 416898 294650 417134
rect 294886 416898 325370 417134
rect 325606 416898 356090 417134
rect 356326 416898 386810 417134
rect 387046 416898 417530 417134
rect 417766 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 64250 399454
rect 64486 399218 94970 399454
rect 95206 399218 125690 399454
rect 125926 399218 156410 399454
rect 156646 399218 187130 399454
rect 187366 399218 217850 399454
rect 218086 399218 248570 399454
rect 248806 399218 279290 399454
rect 279526 399218 310010 399454
rect 310246 399218 340730 399454
rect 340966 399218 371450 399454
rect 371686 399218 402170 399454
rect 402406 399218 432890 399454
rect 433126 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 64250 399134
rect 64486 398898 94970 399134
rect 95206 398898 125690 399134
rect 125926 398898 156410 399134
rect 156646 398898 187130 399134
rect 187366 398898 217850 399134
rect 218086 398898 248570 399134
rect 248806 398898 279290 399134
rect 279526 398898 310010 399134
rect 310246 398898 340730 399134
rect 340966 398898 371450 399134
rect 371686 398898 402170 399134
rect 402406 398898 432890 399134
rect 433126 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect 22564 397578 439644 397620
rect 22564 397342 22606 397578
rect 22842 397342 439366 397578
rect 439602 397342 439644 397578
rect 22564 397300 439644 397342
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect 32132 391458 439644 391500
rect 32132 391222 32174 391458
rect 32410 391222 439366 391458
rect 439602 391222 439644 391458
rect 32132 391180 439644 391222
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 79610 381454
rect 79846 381218 110330 381454
rect 110566 381218 141050 381454
rect 141286 381218 171770 381454
rect 172006 381218 202490 381454
rect 202726 381218 233210 381454
rect 233446 381218 263930 381454
rect 264166 381218 294650 381454
rect 294886 381218 325370 381454
rect 325606 381218 356090 381454
rect 356326 381218 386810 381454
rect 387046 381218 417530 381454
rect 417766 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 79610 381134
rect 79846 380898 110330 381134
rect 110566 380898 141050 381134
rect 141286 380898 171770 381134
rect 172006 380898 202490 381134
rect 202726 380898 233210 381134
rect 233446 380898 263930 381134
rect 264166 380898 294650 381134
rect 294886 380898 325370 381134
rect 325606 380898 356090 381134
rect 356326 380898 386810 381134
rect 387046 380898 417530 381134
rect 417766 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect 60468 371738 500364 371780
rect 60468 371502 60510 371738
rect 60746 371502 500086 371738
rect 500322 371502 500364 371738
rect 60468 371460 500364 371502
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 64250 363454
rect 64486 363218 94970 363454
rect 95206 363218 125690 363454
rect 125926 363218 156410 363454
rect 156646 363218 187130 363454
rect 187366 363218 217850 363454
rect 218086 363218 248570 363454
rect 248806 363218 279290 363454
rect 279526 363218 310010 363454
rect 310246 363218 340730 363454
rect 340966 363218 371450 363454
rect 371686 363218 402170 363454
rect 402406 363218 432890 363454
rect 433126 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 64250 363134
rect 64486 362898 94970 363134
rect 95206 362898 125690 363134
rect 125926 362898 156410 363134
rect 156646 362898 187130 363134
rect 187366 362898 217850 363134
rect 218086 362898 248570 363134
rect 248806 362898 279290 363134
rect 279526 362898 310010 363134
rect 310246 362898 340730 363134
rect 340966 362898 371450 363134
rect 371686 362898 402170 363134
rect 402406 362898 432890 363134
rect 433126 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect 33604 347258 439644 347300
rect 33604 347022 33646 347258
rect 33882 347022 439366 347258
rect 439602 347022 439644 347258
rect 33604 346980 439644 347022
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 79610 345454
rect 79846 345218 110330 345454
rect 110566 345218 141050 345454
rect 141286 345218 171770 345454
rect 172006 345218 202490 345454
rect 202726 345218 233210 345454
rect 233446 345218 263930 345454
rect 264166 345218 294650 345454
rect 294886 345218 325370 345454
rect 325606 345218 356090 345454
rect 356326 345218 386810 345454
rect 387046 345218 417530 345454
rect 417766 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 79610 345134
rect 79846 344898 110330 345134
rect 110566 344898 141050 345134
rect 141286 344898 171770 345134
rect 172006 344898 202490 345134
rect 202726 344898 233210 345134
rect 233446 344898 263930 345134
rect 264166 344898 294650 345134
rect 294886 344898 325370 345134
rect 325606 344898 356090 345134
rect 356326 344898 386810 345134
rect 387046 344898 417530 345134
rect 417766 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect 60468 343858 450684 343900
rect 60468 343622 60510 343858
rect 60746 343622 450406 343858
rect 450642 343622 450684 343858
rect 60468 343580 450684 343622
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 64250 327454
rect 64486 327218 94970 327454
rect 95206 327218 125690 327454
rect 125926 327218 156410 327454
rect 156646 327218 187130 327454
rect 187366 327218 217850 327454
rect 218086 327218 248570 327454
rect 248806 327218 279290 327454
rect 279526 327218 310010 327454
rect 310246 327218 340730 327454
rect 340966 327218 371450 327454
rect 371686 327218 402170 327454
rect 402406 327218 432890 327454
rect 433126 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 64250 327134
rect 64486 326898 94970 327134
rect 95206 326898 125690 327134
rect 125926 326898 156410 327134
rect 156646 326898 187130 327134
rect 187366 326898 217850 327134
rect 218086 326898 248570 327134
rect 248806 326898 279290 327134
rect 279526 326898 310010 327134
rect 310246 326898 340730 327134
rect 340966 326898 371450 327134
rect 371686 326898 402170 327134
rect 402406 326898 432890 327134
rect 433126 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 79610 309454
rect 79846 309218 110330 309454
rect 110566 309218 141050 309454
rect 141286 309218 171770 309454
rect 172006 309218 202490 309454
rect 202726 309218 233210 309454
rect 233446 309218 263930 309454
rect 264166 309218 294650 309454
rect 294886 309218 325370 309454
rect 325606 309218 356090 309454
rect 356326 309218 386810 309454
rect 387046 309218 417530 309454
rect 417766 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 79610 309134
rect 79846 308898 110330 309134
rect 110566 308898 141050 309134
rect 141286 308898 171770 309134
rect 172006 308898 202490 309134
rect 202726 308898 233210 309134
rect 233446 308898 263930 309134
rect 264166 308898 294650 309134
rect 294886 308898 325370 309134
rect 325606 308898 356090 309134
rect 356326 308898 386810 309134
rect 387046 308898 417530 309134
rect 417766 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect 60468 303738 65572 303780
rect 60468 303502 60510 303738
rect 60746 303502 65294 303738
rect 65530 303502 65572 303738
rect 60468 303460 65572 303502
rect 85308 303738 94092 303780
rect 85308 303502 85350 303738
rect 85586 303502 93814 303738
rect 94050 303502 94092 303738
rect 85308 303460 94092 303502
rect 113644 303738 143220 303780
rect 113644 303502 113686 303738
rect 113922 303502 142942 303738
rect 143178 303502 143220 303738
rect 113644 303460 143220 303502
rect 153756 303738 161804 303780
rect 153756 303502 153798 303738
rect 154034 303502 161526 303738
rect 161762 303502 161804 303738
rect 153756 303460 161804 303502
rect 190556 303738 211484 303780
rect 190556 303502 190598 303738
rect 190834 303502 211206 303738
rect 211442 303502 211484 303738
rect 190556 303460 211484 303502
rect 220180 303738 249572 303780
rect 220180 303502 220222 303738
rect 220458 303502 249294 303738
rect 249530 303502 249572 303738
rect 220180 303460 249572 303502
rect 267836 303738 287844 303780
rect 267836 303502 267878 303738
rect 268114 303502 287566 303738
rect 287802 303502 287844 303738
rect 267836 303460 287844 303502
rect 316412 303738 355188 303780
rect 316412 303502 316454 303738
rect 316690 303502 354910 303738
rect 355146 303502 355188 303738
rect 316412 303460 355188 303502
rect 374004 303738 393644 303780
rect 374004 303502 374046 303738
rect 374282 303502 393366 303738
rect 393602 303502 393644 303738
rect 374004 303460 393644 303502
rect 422396 303738 439644 303780
rect 422396 303502 422438 303738
rect 422674 303502 439366 303738
rect 439602 303502 439644 303738
rect 422396 303460 439644 303502
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect 65252 301018 85628 301060
rect 65252 300782 65294 301018
rect 65530 300782 85350 301018
rect 85586 300782 85628 301018
rect 65252 300740 85628 300782
rect 93772 301018 113964 301060
rect 93772 300782 93814 301018
rect 94050 300782 113686 301018
rect 113922 300782 113964 301018
rect 93772 300740 113964 300782
rect 142900 301018 154076 301060
rect 142900 300782 142942 301018
rect 143178 300782 153798 301018
rect 154034 300782 154076 301018
rect 142900 300740 154076 300782
rect 161484 301018 190876 301060
rect 161484 300782 161526 301018
rect 161762 300782 190598 301018
rect 190834 300782 190876 301018
rect 161484 300740 190876 300782
rect 211164 301018 220500 301060
rect 211164 300782 211206 301018
rect 211442 300782 220222 301018
rect 220458 300782 220500 301018
rect 211164 300740 220500 300782
rect 249252 301018 268156 301060
rect 249252 300782 249294 301018
rect 249530 300782 267878 301018
rect 268114 300782 268156 301018
rect 249252 300740 268156 300782
rect 287524 301018 316732 301060
rect 287524 300782 287566 301018
rect 287802 300782 316454 301018
rect 316690 300782 316732 301018
rect 287524 300740 316732 300782
rect 354868 301018 374324 301060
rect 354868 300782 354910 301018
rect 355146 300782 374046 301018
rect 374282 300782 374324 301018
rect 354868 300740 374324 300782
rect 393324 301018 422716 301060
rect 393324 300782 393366 301018
rect 393602 300782 422438 301018
rect 422674 300782 422716 301018
rect 393324 300740 422716 300782
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 64250 291454
rect 64486 291218 94970 291454
rect 95206 291218 125690 291454
rect 125926 291218 156410 291454
rect 156646 291218 187130 291454
rect 187366 291218 217850 291454
rect 218086 291218 248570 291454
rect 248806 291218 279290 291454
rect 279526 291218 310010 291454
rect 310246 291218 340730 291454
rect 340966 291218 371450 291454
rect 371686 291218 402170 291454
rect 402406 291218 432890 291454
rect 433126 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 64250 291134
rect 64486 290898 94970 291134
rect 95206 290898 125690 291134
rect 125926 290898 156410 291134
rect 156646 290898 187130 291134
rect 187366 290898 217850 291134
rect 218086 290898 248570 291134
rect 248806 290898 279290 291134
rect 279526 290898 310010 291134
rect 310246 290898 340730 291134
rect 340966 290898 371450 291134
rect 371686 290898 402170 291134
rect 402406 290898 432890 291134
rect 433126 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect 60468 274498 453444 274540
rect 60468 274262 60510 274498
rect 60746 274262 453166 274498
rect 453402 274262 453444 274498
rect 60468 274220 453444 274262
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 79610 273454
rect 79846 273218 110330 273454
rect 110566 273218 141050 273454
rect 141286 273218 171770 273454
rect 172006 273218 202490 273454
rect 202726 273218 233210 273454
rect 233446 273218 263930 273454
rect 264166 273218 294650 273454
rect 294886 273218 325370 273454
rect 325606 273218 356090 273454
rect 356326 273218 386810 273454
rect 387046 273218 417530 273454
rect 417766 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 79610 273134
rect 79846 272898 110330 273134
rect 110566 272898 141050 273134
rect 141286 272898 171770 273134
rect 172006 272898 202490 273134
rect 202726 272898 233210 273134
rect 233446 272898 263930 273134
rect 264166 272898 294650 273134
rect 294886 272898 325370 273134
rect 325606 272898 356090 273134
rect 356326 272898 386810 273134
rect 387046 272898 417530 273134
rect 417766 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 64250 255454
rect 64486 255218 94970 255454
rect 95206 255218 125690 255454
rect 125926 255218 156410 255454
rect 156646 255218 187130 255454
rect 187366 255218 217850 255454
rect 218086 255218 248570 255454
rect 248806 255218 279290 255454
rect 279526 255218 310010 255454
rect 310246 255218 340730 255454
rect 340966 255218 371450 255454
rect 371686 255218 402170 255454
rect 402406 255218 432890 255454
rect 433126 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 64250 255134
rect 64486 254898 94970 255134
rect 95206 254898 125690 255134
rect 125926 254898 156410 255134
rect 156646 254898 187130 255134
rect 187366 254898 217850 255134
rect 218086 254898 248570 255134
rect 248806 254898 279290 255134
rect 279526 254898 310010 255134
rect 310246 254898 340730 255134
rect 340966 254898 371450 255134
rect 371686 254898 402170 255134
rect 402406 254898 432890 255134
rect 433126 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 79610 237454
rect 79846 237218 110330 237454
rect 110566 237218 141050 237454
rect 141286 237218 171770 237454
rect 172006 237218 202490 237454
rect 202726 237218 233210 237454
rect 233446 237218 263930 237454
rect 264166 237218 294650 237454
rect 294886 237218 325370 237454
rect 325606 237218 356090 237454
rect 356326 237218 386810 237454
rect 387046 237218 417530 237454
rect 417766 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 79610 237134
rect 79846 236898 110330 237134
rect 110566 236898 141050 237134
rect 141286 236898 171770 237134
rect 172006 236898 202490 237134
rect 202726 236898 233210 237134
rect 233446 236898 263930 237134
rect 264166 236898 294650 237134
rect 294886 236898 325370 237134
rect 325606 236898 356090 237134
rect 356326 236898 386810 237134
rect 387046 236898 417530 237134
rect 417766 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 64250 219454
rect 64486 219218 94970 219454
rect 95206 219218 125690 219454
rect 125926 219218 156410 219454
rect 156646 219218 187130 219454
rect 187366 219218 217850 219454
rect 218086 219218 248570 219454
rect 248806 219218 279290 219454
rect 279526 219218 310010 219454
rect 310246 219218 340730 219454
rect 340966 219218 371450 219454
rect 371686 219218 402170 219454
rect 402406 219218 432890 219454
rect 433126 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 64250 219134
rect 64486 218898 94970 219134
rect 95206 218898 125690 219134
rect 125926 218898 156410 219134
rect 156646 218898 187130 219134
rect 187366 218898 217850 219134
rect 218086 218898 248570 219134
rect 248806 218898 279290 219134
rect 279526 218898 310010 219134
rect 310246 218898 340730 219134
rect 340966 218898 371450 219134
rect 371686 218898 402170 219134
rect 402406 218898 432890 219134
rect 433126 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect 60468 213298 468532 213340
rect 60468 213062 60510 213298
rect 60746 213062 468254 213298
rect 468490 213062 468532 213298
rect 60468 213020 468532 213062
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 79610 201454
rect 79846 201218 110330 201454
rect 110566 201218 141050 201454
rect 141286 201218 171770 201454
rect 172006 201218 202490 201454
rect 202726 201218 233210 201454
rect 233446 201218 263930 201454
rect 264166 201218 294650 201454
rect 294886 201218 325370 201454
rect 325606 201218 356090 201454
rect 356326 201218 386810 201454
rect 387046 201218 417530 201454
rect 417766 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 79610 201134
rect 79846 200898 110330 201134
rect 110566 200898 141050 201134
rect 141286 200898 171770 201134
rect 172006 200898 202490 201134
rect 202726 200898 233210 201134
rect 233446 200898 263930 201134
rect 264166 200898 294650 201134
rect 294886 200898 325370 201134
rect 325606 200898 356090 201134
rect 356326 200898 386810 201134
rect 387046 200898 417530 201134
rect 417766 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 64250 183454
rect 64486 183218 94970 183454
rect 95206 183218 125690 183454
rect 125926 183218 156410 183454
rect 156646 183218 187130 183454
rect 187366 183218 217850 183454
rect 218086 183218 248570 183454
rect 248806 183218 279290 183454
rect 279526 183218 310010 183454
rect 310246 183218 340730 183454
rect 340966 183218 371450 183454
rect 371686 183218 402170 183454
rect 402406 183218 432890 183454
rect 433126 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 64250 183134
rect 64486 182898 94970 183134
rect 95206 182898 125690 183134
rect 125926 182898 156410 183134
rect 156646 182898 187130 183134
rect 187366 182898 217850 183134
rect 218086 182898 248570 183134
rect 248806 182898 279290 183134
rect 279526 182898 310010 183134
rect 310246 182898 340730 183134
rect 340966 182898 371450 183134
rect 371686 182898 402170 183134
rect 402406 182898 432890 183134
rect 433126 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect 60468 179298 450684 179340
rect 60468 179062 60510 179298
rect 60746 179062 450406 179298
rect 450642 179062 450684 179298
rect 60468 179020 450684 179062
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 79610 165454
rect 79846 165218 110330 165454
rect 110566 165218 141050 165454
rect 141286 165218 171770 165454
rect 172006 165218 202490 165454
rect 202726 165218 233210 165454
rect 233446 165218 263930 165454
rect 264166 165218 294650 165454
rect 294886 165218 325370 165454
rect 325606 165218 356090 165454
rect 356326 165218 386810 165454
rect 387046 165218 417530 165454
rect 417766 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 79610 165134
rect 79846 164898 110330 165134
rect 110566 164898 141050 165134
rect 141286 164898 171770 165134
rect 172006 164898 202490 165134
rect 202726 164898 233210 165134
rect 233446 164898 263930 165134
rect 264166 164898 294650 165134
rect 294886 164898 325370 165134
rect 325606 164898 356090 165134
rect 356326 164898 386810 165134
rect 387046 164898 417530 165134
rect 417766 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect 60468 160938 471292 160980
rect 60468 160702 60510 160938
rect 60746 160702 471014 160938
rect 471250 160702 471292 160938
rect 60468 160660 471292 160702
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 125690 147454
rect 125926 147218 156410 147454
rect 156646 147218 187130 147454
rect 187366 147218 217850 147454
rect 218086 147218 248570 147454
rect 248806 147218 279290 147454
rect 279526 147218 310010 147454
rect 310246 147218 340730 147454
rect 340966 147218 371450 147454
rect 371686 147218 402170 147454
rect 402406 147218 432890 147454
rect 433126 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 125690 147134
rect 125926 146898 156410 147134
rect 156646 146898 187130 147134
rect 187366 146898 217850 147134
rect 218086 146898 248570 147134
rect 248806 146898 279290 147134
rect 279526 146898 310010 147134
rect 310246 146898 340730 147134
rect 340966 146898 371450 147134
rect 371686 146898 402170 147134
rect 402406 146898 432890 147134
rect 433126 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 79610 129454
rect 79846 129218 110330 129454
rect 110566 129218 141050 129454
rect 141286 129218 171770 129454
rect 172006 129218 202490 129454
rect 202726 129218 233210 129454
rect 233446 129218 263930 129454
rect 264166 129218 294650 129454
rect 294886 129218 325370 129454
rect 325606 129218 356090 129454
rect 356326 129218 386810 129454
rect 387046 129218 417530 129454
rect 417766 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 79610 129134
rect 79846 128898 110330 129134
rect 110566 128898 141050 129134
rect 141286 128898 171770 129134
rect 172006 128898 202490 129134
rect 202726 128898 233210 129134
rect 233446 128898 263930 129134
rect 264166 128898 294650 129134
rect 294886 128898 325370 129134
rect 325606 128898 356090 129134
rect 356326 128898 386810 129134
rect 387046 128898 417530 129134
rect 417766 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 64250 111454
rect 64486 111218 94970 111454
rect 95206 111218 125690 111454
rect 125926 111218 156410 111454
rect 156646 111218 187130 111454
rect 187366 111218 217850 111454
rect 218086 111218 248570 111454
rect 248806 111218 279290 111454
rect 279526 111218 310010 111454
rect 310246 111218 340730 111454
rect 340966 111218 371450 111454
rect 371686 111218 402170 111454
rect 402406 111218 432890 111454
rect 433126 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 64250 111134
rect 64486 110898 94970 111134
rect 95206 110898 125690 111134
rect 125926 110898 156410 111134
rect 156646 110898 187130 111134
rect 187366 110898 217850 111134
rect 218086 110898 248570 111134
rect 248806 110898 279290 111134
rect 279526 110898 310010 111134
rect 310246 110898 340730 111134
rect 340966 110898 371450 111134
rect 371686 110898 402170 111134
rect 402406 110898 432890 111134
rect 433126 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 79610 93454
rect 79846 93218 110330 93454
rect 110566 93218 141050 93454
rect 141286 93218 171770 93454
rect 172006 93218 202490 93454
rect 202726 93218 233210 93454
rect 233446 93218 263930 93454
rect 264166 93218 294650 93454
rect 294886 93218 325370 93454
rect 325606 93218 356090 93454
rect 356326 93218 386810 93454
rect 387046 93218 417530 93454
rect 417766 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 79610 93134
rect 79846 92898 110330 93134
rect 110566 92898 141050 93134
rect 141286 92898 171770 93134
rect 172006 92898 202490 93134
rect 202726 92898 233210 93134
rect 233446 92898 263930 93134
rect 264166 92898 294650 93134
rect 294886 92898 325370 93134
rect 325606 92898 356090 93134
rect 356326 92898 386810 93134
rect 387046 92898 417530 93134
rect 417766 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 64250 75454
rect 64486 75218 94970 75454
rect 95206 75218 125690 75454
rect 125926 75218 156410 75454
rect 156646 75218 187130 75454
rect 187366 75218 217850 75454
rect 218086 75218 248570 75454
rect 248806 75218 279290 75454
rect 279526 75218 310010 75454
rect 310246 75218 340730 75454
rect 340966 75218 371450 75454
rect 371686 75218 402170 75454
rect 402406 75218 432890 75454
rect 433126 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 64250 75134
rect 64486 74898 94970 75134
rect 95206 74898 125690 75134
rect 125926 74898 156410 75134
rect 156646 74898 187130 75134
rect 187366 74898 217850 75134
rect 218086 74898 248570 75134
rect 248806 74898 279290 75134
rect 279526 74898 310010 75134
rect 310246 74898 340730 75134
rect 340966 74898 371450 75134
rect 371686 74898 402170 75134
rect 402406 74898 432890 75134
rect 433126 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect 61940 4538 309372 4580
rect 61940 4302 61982 4538
rect 62218 4302 309094 4538
rect 309330 4302 309372 4538
rect 61940 4260 309372 4302
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj_systollic  mprj
timestamp 1667209117
transform 1 0 60000 0 1 60000
box 0 0 380000 480000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 542000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 542000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 542000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 542000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 542000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 542000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 542000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 542000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 542000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 542000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 542000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 542000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 542000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 542000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 542000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 542000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 542000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 542000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 542000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 542000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 542000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 542000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 542000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 542000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 542000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 542000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 542000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 542000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 542000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 542000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 542000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 542000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 542000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 542000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 542000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 542000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 542000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 542000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 542000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 542000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 542000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 542000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 542000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 542000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 542000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 542000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 542000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 542000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 542000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 542000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 542000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 542000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 542000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 542000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 542000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 542000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 542000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 542000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 542000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 542000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 542000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 542000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 542000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 542000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 542000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 542000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 542000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 542000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 542000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 542000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 542000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 542000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 542000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 542000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 542000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 542000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 542000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 542000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 542000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 542000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 542000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 542000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 542000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 542000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 542000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 542000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
