VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_systollic
  CLASS BLOCK ;
  FOREIGN user_proj_systollic ;
  ORIGIN 0.000 0.000 ;
  SIZE 1900.000 BY 2400.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 156.440 1900.000 157.040 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1186.640 1900.000 1187.240 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 2396.000 489.810 2400.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1652.440 1900.000 1653.040 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 2396.000 380.330 2400.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2305.240 1900.000 2305.840 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 2396.000 557.430 2400.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 2396.000 309.490 2400.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 2396.000 418.970 2400.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1839.440 1900.000 1840.040 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2247.440 4.000 2248.040 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 2396.000 1108.050 2400.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 2396.000 351.350 2400.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 2396.000 737.750 2400.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1798.640 4.000 1799.240 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 2396.000 1217.530 2400.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.170 2396.000 1011.450 2400.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1666.040 1900.000 1666.640 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 40.840 1900.000 41.440 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.750 2396.000 1781.030 2400.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 489.640 1900.000 490.240 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1506.240 1900.000 1506.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 2396.000 792.490 2400.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.240 4.000 1421.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 996.240 1900.000 996.840 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 955.440 1900.000 956.040 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 2396.000 1040.430 2400.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 2396.000 515.570 2400.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.130 0.000 1552.410 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 2396.000 145.270 2400.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1013.240 1900.000 1013.840 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2176.040 4.000 2176.640 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2220.240 4.000 2220.840 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 0.000 1413.950 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 2396.000 158.150 2400.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.130 2396.000 1230.410 2400.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1115.240 1900.000 1115.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2376.640 1900.000 2377.240 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 2396.000 22.910 2400.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 2396.000 1066.190 2400.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1825.840 1900.000 1826.440 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2101.240 1900.000 2101.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.190 0.000 1304.470 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.840 4.000 1928.440 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 2396.000 48.670 2400.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2264.440 4.000 2265.040 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 2396.000 174.250 2400.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1608.240 4.000 1608.840 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 2396.000 1397.850 2400.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 2396.000 1301.250 2400.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.610 2396.000 1822.890 2400.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1550.440 4.000 1551.040 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2393.640 4.000 2394.240 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2145.440 4.000 2146.040 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1767.870 2396.000 1768.150 2400.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2247.440 1900.000 2248.040 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1910.840 1900.000 1911.440 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 720.840 1900.000 721.440 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1635.440 1900.000 1636.040 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2172.640 1900.000 2173.240 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1927.840 1900.000 1928.440 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 0.000 1607.150 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2118.240 4.000 2118.840 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 98.640 1900.000 99.240 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 459.040 1900.000 459.640 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1492.640 4.000 1493.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 2396.000 200.010 2400.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 214.240 1900.000 214.840 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1434.840 1900.000 1435.440 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 2396.000 1810.010 2400.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2145.440 1900.000 2146.040 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.670 0.000 1896.950 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1870.040 1900.000 1870.640 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.350 2396.000 1877.630 2400.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1693.240 1900.000 1693.840 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 2396.000 187.130 2400.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.790 0.000 1884.070 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 431.840 1900.000 432.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1577.640 1900.000 1578.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 2396.000 847.230 2400.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 2396.000 641.150 2400.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2131.840 4.000 2132.440 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1098.240 1900.000 1098.840 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 2396.000 1452.590 2400.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1332.840 1900.000 1333.440 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 836.440 1900.000 837.040 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 2396.000 708.770 2400.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 2396.000 119.510 2400.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2216.840 1900.000 2217.440 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1652.440 4.000 1653.040 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1594.640 1900.000 1595.240 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 445.440 1900.000 446.040 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 2396.000 927.730 2400.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 795.640 1900.000 796.240 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 2396.000 1285.150 2400.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1696.640 4.000 1697.240 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1608.240 1900.000 1608.840 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 561.040 1900.000 561.640 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 2396.000 1343.110 2400.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 2396.000 628.270 2400.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 2396.000 1478.350 2400.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1533.440 1900.000 1534.040 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1581.040 4.000 1581.640 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 2396.000 1204.650 2400.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 139.440 1900.000 140.040 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2278.040 4.000 2278.640 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 241.440 1900.000 242.040 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2366.440 4.000 2367.040 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.990 0.000 1594.270 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 0.000 1855.090 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1795.240 1900.000 1795.840 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1142.440 1900.000 1143.040 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2057.040 1900.000 2057.640 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 2396.000 1381.750 2400.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2206.640 4.000 2207.240 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1373.640 1900.000 1374.240 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 649.440 1900.000 650.040 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.840 4.000 1452.440 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1972.040 1900.000 1972.640 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1519.840 1900.000 1520.440 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 0.000 1661.890 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 68.040 1900.000 68.640 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 2396.000 544.550 2400.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 0.000 1523.430 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 2396.000 750.630 2400.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1829.240 4.000 1829.840 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 2396.000 1436.490 2400.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 2396.000 1835.770 2400.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1173.040 1900.000 1173.640 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1213.840 1900.000 1214.440 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1897.240 1900.000 1897.840 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 2396.000 476.930 2400.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1203.640 4.000 1204.240 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 0.000 1401.070 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 2396.000 1272.270 2400.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2189.640 4.000 2190.240 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.630 2396.000 1793.910 2400.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 635.840 1900.000 636.440 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 2396.000 1533.090 2400.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 0.000 1826.110 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2335.840 4.000 2336.440 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 751.440 1900.000 752.040 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2274.640 1900.000 2275.240 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2060.440 4.000 2061.040 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 2396.000 654.030 2400.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1812.240 1900.000 1812.840 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1084.640 1900.000 1085.240 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 765.040 1900.000 765.640 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 618.840 1900.000 619.440 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 2396.000 296.610 2400.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 183.640 1900.000 184.240 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1621.840 1900.000 1622.440 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1955.040 1900.000 1955.640 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 822.840 1900.000 823.440 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 897.640 1900.000 898.240 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.350 0.000 1716.630 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 911.240 1900.000 911.840 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.910 2396.000 1549.190 2400.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 2396.000 612.170 2400.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1768.040 1900.000 1768.640 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 2396.000 502.690 2400.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 2396.000 267.630 2400.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 2396.000 998.570 2400.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2233.840 4.000 2234.440 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 258.440 1900.000 259.040 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 401.240 1900.000 401.840 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1914.240 4.000 1914.840 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1244.440 1900.000 1245.040 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1479.040 4.000 1479.640 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 2396.000 1739.170 2400.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1900.640 4.000 1901.240 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1026.840 1900.000 1027.440 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1404.240 1900.000 1404.840 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 2396.000 254.750 2400.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 0.000 1375.310 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1740.840 4.000 1741.440 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 2396.000 872.990 2400.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 2396.000 1053.310 2400.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 2396.000 1327.010 2400.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 2396.000 1700.530 2400.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 2396.000 666.910 2400.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2131.840 1900.000 2132.440 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 707.240 1900.000 707.840 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 285.640 1900.000 286.240 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 2396.000 132.390 2400.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 2396.000 1726.290 2400.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1754.440 4.000 1755.040 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 10.240 1900.000 10.840 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2159.040 1900.000 2159.640 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1200.240 1900.000 1200.840 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1302.240 1900.000 1302.840 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 170.040 1900.000 170.640 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2349.440 4.000 2350.040 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 591.640 1900.000 592.240 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2322.240 4.000 2322.840 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2332.440 1900.000 2333.040 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 2396.000 1162.790 2400.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1040.440 1900.000 1041.040 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 2396.000 956.710 2400.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1230.840 1900.000 1231.440 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2029.840 4.000 2030.440 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 533.840 1900.000 534.440 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 2396.000 228.990 2400.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 2396.000 985.690 2400.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 125.840 1900.000 126.440 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 2396.000 1645.790 2400.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.840 4.000 1639.440 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 2396.000 1465.470 2400.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 809.240 1900.000 809.840 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 2396.000 586.410 2400.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 2396.000 435.070 2400.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 2396.000 364.230 2400.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 272.040 1900.000 272.640 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.470 2396.000 1864.750 2400.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 2396.000 531.670 2400.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1247.840 4.000 1248.440 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1669.440 4.000 1670.040 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1315.840 1900.000 1316.440 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1258.040 1900.000 1258.640 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.990 2396.000 1755.270 2400.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 2396.000 1410.730 2400.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 2396.000 805.370 2400.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.730 0.000 1649.010 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1870.040 4.000 1870.640 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1390.640 1900.000 1391.240 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 693.640 1900.000 694.240 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 503.240 1900.000 503.840 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 0.000 1484.790 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.150 2396.000 1684.430 2400.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 2396.000 599.290 2400.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2074.040 4.000 2074.640 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 2396.000 834.350 2400.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 418.240 1900.000 418.840 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 81.640 1900.000 82.240 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 676.640 1900.000 677.240 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 578.040 1900.000 578.640 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2016.240 4.000 2016.840 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 2396.000 241.870 2400.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 0.000 1703.750 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 2396.000 90.530 2400.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 200.640 1900.000 201.240 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1346.440 1900.000 1347.040 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 2396.000 943.830 2400.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 2396.000 889.090 2400.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 2396.000 901.970 2400.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 0.000 1581.390 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.090 0.000 1771.370 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 2396.000 1574.950 2400.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 2396.000 460.830 2400.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 2396.000 683.010 2400.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.850 0.000 1636.130 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2380.040 4.000 2380.640 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 2396.000 1520.210 2400.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 227.840 1900.000 228.440 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2363.040 1900.000 2363.640 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1842.840 4.000 1843.440 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.790 2396.000 1562.070 2400.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1475.640 1900.000 1476.240 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 2396.000 763.510 2400.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.590 2396.000 1851.870 2400.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1448.440 1900.000 1449.040 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 2396.000 1175.670 2400.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 2396.000 1423.610 2400.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1883.640 1900.000 1884.240 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 0.000 1539.530 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.840 4.000 1146.440 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 2396.000 1024.330 2400.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2288.240 1900.000 2288.840 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1071.040 1900.000 1071.640 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1462.040 1900.000 1462.640 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 0.000 1346.330 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1594.640 4.000 1595.240 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2029.840 1900.000 2030.440 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.450 0.000 1732.730 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 778.640 1900.000 779.240 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1723.840 1900.000 1724.440 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 605.240 1900.000 605.840 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 547.440 1900.000 548.040 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2261.040 1900.000 2261.640 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1128.840 1900.000 1129.440 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.410 2396.000 1629.690 2400.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1417.840 1900.000 1418.440 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 2396.000 1890.510 2400.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 2396.000 1658.670 2400.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 2396.000 393.210 2400.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 2396.000 35.790 2400.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 924.840 1900.000 925.440 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1492.640 1900.000 1493.240 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.750 0.000 1620.030 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1999.240 1900.000 1999.840 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1465.440 4.000 1466.040 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 2396.000 1713.410 2400.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1887.040 4.000 1887.640 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 54.440 1900.000 55.040 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2291.640 4.000 2292.240 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1856.440 4.000 1857.040 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 360.440 1900.000 361.040 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 112.240 1900.000 112.840 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 880.640 1900.000 881.240 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2012.840 1900.000 2013.440 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 2396.000 776.390 2400.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 2396.000 447.950 2400.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2230.440 1900.000 2231.040 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.240 4.000 1625.840 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 2396.000 325.590 2400.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1985.640 1900.000 1986.240 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.110 2396.000 1259.390 2400.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2046.840 4.000 2047.440 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 2396.000 1494.450 2400.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 2396.000 1603.930 2400.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.530 2396.000 1616.810 2400.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 2396.000 914.850 2400.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.690 0.000 1867.970 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 663.040 1900.000 663.640 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2104.640 4.000 2105.240 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 2396.000 860.110 2400.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 23.840 1900.000 24.440 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1785.040 4.000 1785.640 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1737.440 1900.000 1738.040 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2203.240 1900.000 2203.840 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1292.040 4.000 1292.640 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1567.440 4.000 1568.040 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 476.040 1900.000 476.640 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2087.640 1900.000 2088.240 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 2396.000 570.310 2400.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1781.640 1900.000 1782.240 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.070 0.000 1800.350 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 737.840 1900.000 738.440 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 2396.000 406.090 2400.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 299.240 1900.000 299.840 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1989.040 4.000 1989.640 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.070 0.000 1317.350 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2070.640 1900.000 2071.240 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 329.840 1900.000 330.440 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2162.440 4.000 2163.040 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 2396.000 1095.170 2400.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2087.640 4.000 2088.240 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2305.240 4.000 2305.840 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2388.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2388.400 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 867.040 1900.000 867.640 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1958.440 4.000 1959.040 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 2396.000 695.890 2400.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 2396.000 212.890 2400.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1683.040 4.000 1683.640 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1305.640 4.000 1306.240 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2189.640 1900.000 2190.240 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2043.440 1900.000 2044.040 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1156.040 1900.000 1156.640 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 316.240 1900.000 316.840 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 2396.000 721.650 2400.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 2396.000 1368.870 2400.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 0.000 1842.210 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 938.440 1900.000 939.040 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1944.840 4.000 1945.440 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 2396.000 77.650 2400.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1751.040 1900.000 1751.640 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 2396.000 1671.550 2400.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 2396.000 1120.930 2400.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1360.040 1900.000 1360.640 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.330 0.000 1745.610 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 2396.000 1079.070 2400.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 0.000 1674.770 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 343.440 1900.000 344.040 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 982.640 1900.000 983.240 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 2396.000 103.410 2400.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2390.240 1900.000 2390.840 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1550.440 1900.000 1551.040 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 2396.000 969.590 2400.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 2396.000 1507.330 2400.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1972.040 4.000 1972.640 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1710.240 1900.000 1710.840 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.550 2396.000 1587.830 2400.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2114.840 1900.000 2115.440 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1057.440 1900.000 1058.040 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 2396.000 1355.990 2400.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 2396.000 61.550 2400.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1679.640 1900.000 1680.240 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 969.040 1900.000 969.640 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 374.040 1900.000 374.640 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1275.040 1900.000 1275.640 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 2396.000 1314.130 2400.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2318.840 1900.000 2319.440 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 387.640 1900.000 388.240 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1564.040 1900.000 1564.640 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 2349.440 1900.000 2350.040 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 2396.000 1246.510 2400.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 520.240 1900.000 520.840 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 0.000 1442.930 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.590 0.000 1690.870 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.040 4.000 1768.640 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 2396.000 283.730 2400.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 2396.000 818.250 2400.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 2396.000 338.470 2400.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 2396.000 1191.770 2400.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 853.440 1900.000 854.040 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1363.440 4.000 1364.040 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1941.440 1900.000 1942.040 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1853.040 1900.000 1853.640 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.430 0.000 1278.710 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 2396.000 1149.910 2400.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 2396.000 1137.030 2400.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2002.640 4.000 2003.240 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 2396.000 6.810 2400.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1812.240 4.000 1812.840 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1896.000 1288.640 1900.000 1289.240 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1894.280 2388.245 ;
      LAYER met1 ;
        RECT 0.070 9.220 1896.970 2388.400 ;
      LAYER met2 ;
        RECT 0.100 2395.720 6.250 2396.730 ;
        RECT 7.090 2395.720 22.350 2396.730 ;
        RECT 23.190 2395.720 35.230 2396.730 ;
        RECT 36.070 2395.720 48.110 2396.730 ;
        RECT 48.950 2395.720 60.990 2396.730 ;
        RECT 61.830 2395.720 77.090 2396.730 ;
        RECT 77.930 2395.720 89.970 2396.730 ;
        RECT 90.810 2395.720 102.850 2396.730 ;
        RECT 103.690 2395.720 118.950 2396.730 ;
        RECT 119.790 2395.720 131.830 2396.730 ;
        RECT 132.670 2395.720 144.710 2396.730 ;
        RECT 145.550 2395.720 157.590 2396.730 ;
        RECT 158.430 2395.720 173.690 2396.730 ;
        RECT 174.530 2395.720 186.570 2396.730 ;
        RECT 187.410 2395.720 199.450 2396.730 ;
        RECT 200.290 2395.720 212.330 2396.730 ;
        RECT 213.170 2395.720 228.430 2396.730 ;
        RECT 229.270 2395.720 241.310 2396.730 ;
        RECT 242.150 2395.720 254.190 2396.730 ;
        RECT 255.030 2395.720 267.070 2396.730 ;
        RECT 267.910 2395.720 283.170 2396.730 ;
        RECT 284.010 2395.720 296.050 2396.730 ;
        RECT 296.890 2395.720 308.930 2396.730 ;
        RECT 309.770 2395.720 325.030 2396.730 ;
        RECT 325.870 2395.720 337.910 2396.730 ;
        RECT 338.750 2395.720 350.790 2396.730 ;
        RECT 351.630 2395.720 363.670 2396.730 ;
        RECT 364.510 2395.720 379.770 2396.730 ;
        RECT 380.610 2395.720 392.650 2396.730 ;
        RECT 393.490 2395.720 405.530 2396.730 ;
        RECT 406.370 2395.720 418.410 2396.730 ;
        RECT 419.250 2395.720 434.510 2396.730 ;
        RECT 435.350 2395.720 447.390 2396.730 ;
        RECT 448.230 2395.720 460.270 2396.730 ;
        RECT 461.110 2395.720 476.370 2396.730 ;
        RECT 477.210 2395.720 489.250 2396.730 ;
        RECT 490.090 2395.720 502.130 2396.730 ;
        RECT 502.970 2395.720 515.010 2396.730 ;
        RECT 515.850 2395.720 531.110 2396.730 ;
        RECT 531.950 2395.720 543.990 2396.730 ;
        RECT 544.830 2395.720 556.870 2396.730 ;
        RECT 557.710 2395.720 569.750 2396.730 ;
        RECT 570.590 2395.720 585.850 2396.730 ;
        RECT 586.690 2395.720 598.730 2396.730 ;
        RECT 599.570 2395.720 611.610 2396.730 ;
        RECT 612.450 2395.720 627.710 2396.730 ;
        RECT 628.550 2395.720 640.590 2396.730 ;
        RECT 641.430 2395.720 653.470 2396.730 ;
        RECT 654.310 2395.720 666.350 2396.730 ;
        RECT 667.190 2395.720 682.450 2396.730 ;
        RECT 683.290 2395.720 695.330 2396.730 ;
        RECT 696.170 2395.720 708.210 2396.730 ;
        RECT 709.050 2395.720 721.090 2396.730 ;
        RECT 721.930 2395.720 737.190 2396.730 ;
        RECT 738.030 2395.720 750.070 2396.730 ;
        RECT 750.910 2395.720 762.950 2396.730 ;
        RECT 763.790 2395.720 775.830 2396.730 ;
        RECT 776.670 2395.720 791.930 2396.730 ;
        RECT 792.770 2395.720 804.810 2396.730 ;
        RECT 805.650 2395.720 817.690 2396.730 ;
        RECT 818.530 2395.720 833.790 2396.730 ;
        RECT 834.630 2395.720 846.670 2396.730 ;
        RECT 847.510 2395.720 859.550 2396.730 ;
        RECT 860.390 2395.720 872.430 2396.730 ;
        RECT 873.270 2395.720 888.530 2396.730 ;
        RECT 889.370 2395.720 901.410 2396.730 ;
        RECT 902.250 2395.720 914.290 2396.730 ;
        RECT 915.130 2395.720 927.170 2396.730 ;
        RECT 928.010 2395.720 943.270 2396.730 ;
        RECT 944.110 2395.720 956.150 2396.730 ;
        RECT 956.990 2395.720 969.030 2396.730 ;
        RECT 969.870 2395.720 985.130 2396.730 ;
        RECT 985.970 2395.720 998.010 2396.730 ;
        RECT 998.850 2395.720 1010.890 2396.730 ;
        RECT 1011.730 2395.720 1023.770 2396.730 ;
        RECT 1024.610 2395.720 1039.870 2396.730 ;
        RECT 1040.710 2395.720 1052.750 2396.730 ;
        RECT 1053.590 2395.720 1065.630 2396.730 ;
        RECT 1066.470 2395.720 1078.510 2396.730 ;
        RECT 1079.350 2395.720 1094.610 2396.730 ;
        RECT 1095.450 2395.720 1107.490 2396.730 ;
        RECT 1108.330 2395.720 1120.370 2396.730 ;
        RECT 1121.210 2395.720 1136.470 2396.730 ;
        RECT 1137.310 2395.720 1149.350 2396.730 ;
        RECT 1150.190 2395.720 1162.230 2396.730 ;
        RECT 1163.070 2395.720 1175.110 2396.730 ;
        RECT 1175.950 2395.720 1191.210 2396.730 ;
        RECT 1192.050 2395.720 1204.090 2396.730 ;
        RECT 1204.930 2395.720 1216.970 2396.730 ;
        RECT 1217.810 2395.720 1229.850 2396.730 ;
        RECT 1230.690 2395.720 1245.950 2396.730 ;
        RECT 1246.790 2395.720 1258.830 2396.730 ;
        RECT 1259.670 2395.720 1271.710 2396.730 ;
        RECT 1272.550 2395.720 1284.590 2396.730 ;
        RECT 1285.430 2395.720 1300.690 2396.730 ;
        RECT 1301.530 2395.720 1313.570 2396.730 ;
        RECT 1314.410 2395.720 1326.450 2396.730 ;
        RECT 1327.290 2395.720 1342.550 2396.730 ;
        RECT 1343.390 2395.720 1355.430 2396.730 ;
        RECT 1356.270 2395.720 1368.310 2396.730 ;
        RECT 1369.150 2395.720 1381.190 2396.730 ;
        RECT 1382.030 2395.720 1397.290 2396.730 ;
        RECT 1398.130 2395.720 1410.170 2396.730 ;
        RECT 1411.010 2395.720 1423.050 2396.730 ;
        RECT 1423.890 2395.720 1435.930 2396.730 ;
        RECT 1436.770 2395.720 1452.030 2396.730 ;
        RECT 1452.870 2395.720 1464.910 2396.730 ;
        RECT 1465.750 2395.720 1477.790 2396.730 ;
        RECT 1478.630 2395.720 1493.890 2396.730 ;
        RECT 1494.730 2395.720 1506.770 2396.730 ;
        RECT 1507.610 2395.720 1519.650 2396.730 ;
        RECT 1520.490 2395.720 1532.530 2396.730 ;
        RECT 1533.370 2395.720 1548.630 2396.730 ;
        RECT 1549.470 2395.720 1561.510 2396.730 ;
        RECT 1562.350 2395.720 1574.390 2396.730 ;
        RECT 1575.230 2395.720 1587.270 2396.730 ;
        RECT 1588.110 2395.720 1603.370 2396.730 ;
        RECT 1604.210 2395.720 1616.250 2396.730 ;
        RECT 1617.090 2395.720 1629.130 2396.730 ;
        RECT 1629.970 2395.720 1645.230 2396.730 ;
        RECT 1646.070 2395.720 1658.110 2396.730 ;
        RECT 1658.950 2395.720 1670.990 2396.730 ;
        RECT 1671.830 2395.720 1683.870 2396.730 ;
        RECT 1684.710 2395.720 1699.970 2396.730 ;
        RECT 1700.810 2395.720 1712.850 2396.730 ;
        RECT 1713.690 2395.720 1725.730 2396.730 ;
        RECT 1726.570 2395.720 1738.610 2396.730 ;
        RECT 1739.450 2395.720 1754.710 2396.730 ;
        RECT 1755.550 2395.720 1767.590 2396.730 ;
        RECT 1768.430 2395.720 1780.470 2396.730 ;
        RECT 1781.310 2395.720 1793.350 2396.730 ;
        RECT 1794.190 2395.720 1809.450 2396.730 ;
        RECT 1810.290 2395.720 1822.330 2396.730 ;
        RECT 1823.170 2395.720 1835.210 2396.730 ;
        RECT 1836.050 2395.720 1851.310 2396.730 ;
        RECT 1852.150 2395.720 1864.190 2396.730 ;
        RECT 1865.030 2395.720 1877.070 2396.730 ;
        RECT 1877.910 2395.720 1889.950 2396.730 ;
        RECT 1890.790 2395.720 1896.940 2396.730 ;
        RECT 0.100 4.280 1896.940 2395.720 ;
        RECT 0.650 4.000 12.690 4.280 ;
        RECT 13.530 4.000 25.570 4.280 ;
        RECT 26.410 4.000 38.450 4.280 ;
        RECT 39.290 4.000 54.550 4.280 ;
        RECT 55.390 4.000 67.430 4.280 ;
        RECT 68.270 4.000 80.310 4.280 ;
        RECT 81.150 4.000 93.190 4.280 ;
        RECT 94.030 4.000 109.290 4.280 ;
        RECT 110.130 4.000 122.170 4.280 ;
        RECT 123.010 4.000 135.050 4.280 ;
        RECT 135.890 4.000 147.930 4.280 ;
        RECT 148.770 4.000 164.030 4.280 ;
        RECT 164.870 4.000 176.910 4.280 ;
        RECT 177.750 4.000 189.790 4.280 ;
        RECT 190.630 4.000 205.890 4.280 ;
        RECT 206.730 4.000 218.770 4.280 ;
        RECT 219.610 4.000 231.650 4.280 ;
        RECT 232.490 4.000 244.530 4.280 ;
        RECT 245.370 4.000 260.630 4.280 ;
        RECT 261.470 4.000 273.510 4.280 ;
        RECT 274.350 4.000 286.390 4.280 ;
        RECT 287.230 4.000 299.270 4.280 ;
        RECT 300.110 4.000 315.370 4.280 ;
        RECT 316.210 4.000 328.250 4.280 ;
        RECT 329.090 4.000 341.130 4.280 ;
        RECT 341.970 4.000 357.230 4.280 ;
        RECT 358.070 4.000 370.110 4.280 ;
        RECT 370.950 4.000 382.990 4.280 ;
        RECT 383.830 4.000 395.870 4.280 ;
        RECT 396.710 4.000 411.970 4.280 ;
        RECT 412.810 4.000 424.850 4.280 ;
        RECT 425.690 4.000 437.730 4.280 ;
        RECT 438.570 4.000 450.610 4.280 ;
        RECT 451.450 4.000 466.710 4.280 ;
        RECT 467.550 4.000 479.590 4.280 ;
        RECT 480.430 4.000 492.470 4.280 ;
        RECT 493.310 4.000 505.350 4.280 ;
        RECT 506.190 4.000 521.450 4.280 ;
        RECT 522.290 4.000 534.330 4.280 ;
        RECT 535.170 4.000 547.210 4.280 ;
        RECT 548.050 4.000 563.310 4.280 ;
        RECT 564.150 4.000 576.190 4.280 ;
        RECT 577.030 4.000 589.070 4.280 ;
        RECT 589.910 4.000 601.950 4.280 ;
        RECT 602.790 4.000 618.050 4.280 ;
        RECT 618.890 4.000 630.930 4.280 ;
        RECT 631.770 4.000 643.810 4.280 ;
        RECT 644.650 4.000 656.690 4.280 ;
        RECT 657.530 4.000 672.790 4.280 ;
        RECT 673.630 4.000 685.670 4.280 ;
        RECT 686.510 4.000 698.550 4.280 ;
        RECT 699.390 4.000 714.650 4.280 ;
        RECT 715.490 4.000 727.530 4.280 ;
        RECT 728.370 4.000 740.410 4.280 ;
        RECT 741.250 4.000 753.290 4.280 ;
        RECT 754.130 4.000 769.390 4.280 ;
        RECT 770.230 4.000 782.270 4.280 ;
        RECT 783.110 4.000 795.150 4.280 ;
        RECT 795.990 4.000 808.030 4.280 ;
        RECT 808.870 4.000 824.130 4.280 ;
        RECT 824.970 4.000 837.010 4.280 ;
        RECT 837.850 4.000 849.890 4.280 ;
        RECT 850.730 4.000 865.990 4.280 ;
        RECT 866.830 4.000 878.870 4.280 ;
        RECT 879.710 4.000 891.750 4.280 ;
        RECT 892.590 4.000 904.630 4.280 ;
        RECT 905.470 4.000 920.730 4.280 ;
        RECT 921.570 4.000 933.610 4.280 ;
        RECT 934.450 4.000 946.490 4.280 ;
        RECT 947.330 4.000 959.370 4.280 ;
        RECT 960.210 4.000 975.470 4.280 ;
        RECT 976.310 4.000 988.350 4.280 ;
        RECT 989.190 4.000 1001.230 4.280 ;
        RECT 1002.070 4.000 1014.110 4.280 ;
        RECT 1014.950 4.000 1030.210 4.280 ;
        RECT 1031.050 4.000 1043.090 4.280 ;
        RECT 1043.930 4.000 1055.970 4.280 ;
        RECT 1056.810 4.000 1072.070 4.280 ;
        RECT 1072.910 4.000 1084.950 4.280 ;
        RECT 1085.790 4.000 1097.830 4.280 ;
        RECT 1098.670 4.000 1110.710 4.280 ;
        RECT 1111.550 4.000 1126.810 4.280 ;
        RECT 1127.650 4.000 1139.690 4.280 ;
        RECT 1140.530 4.000 1152.570 4.280 ;
        RECT 1153.410 4.000 1165.450 4.280 ;
        RECT 1166.290 4.000 1181.550 4.280 ;
        RECT 1182.390 4.000 1194.430 4.280 ;
        RECT 1195.270 4.000 1207.310 4.280 ;
        RECT 1208.150 4.000 1223.410 4.280 ;
        RECT 1224.250 4.000 1236.290 4.280 ;
        RECT 1237.130 4.000 1249.170 4.280 ;
        RECT 1250.010 4.000 1262.050 4.280 ;
        RECT 1262.890 4.000 1278.150 4.280 ;
        RECT 1278.990 4.000 1291.030 4.280 ;
        RECT 1291.870 4.000 1303.910 4.280 ;
        RECT 1304.750 4.000 1316.790 4.280 ;
        RECT 1317.630 4.000 1332.890 4.280 ;
        RECT 1333.730 4.000 1345.770 4.280 ;
        RECT 1346.610 4.000 1358.650 4.280 ;
        RECT 1359.490 4.000 1374.750 4.280 ;
        RECT 1375.590 4.000 1387.630 4.280 ;
        RECT 1388.470 4.000 1400.510 4.280 ;
        RECT 1401.350 4.000 1413.390 4.280 ;
        RECT 1414.230 4.000 1429.490 4.280 ;
        RECT 1430.330 4.000 1442.370 4.280 ;
        RECT 1443.210 4.000 1455.250 4.280 ;
        RECT 1456.090 4.000 1468.130 4.280 ;
        RECT 1468.970 4.000 1484.230 4.280 ;
        RECT 1485.070 4.000 1497.110 4.280 ;
        RECT 1497.950 4.000 1509.990 4.280 ;
        RECT 1510.830 4.000 1522.870 4.280 ;
        RECT 1523.710 4.000 1538.970 4.280 ;
        RECT 1539.810 4.000 1551.850 4.280 ;
        RECT 1552.690 4.000 1564.730 4.280 ;
        RECT 1565.570 4.000 1580.830 4.280 ;
        RECT 1581.670 4.000 1593.710 4.280 ;
        RECT 1594.550 4.000 1606.590 4.280 ;
        RECT 1607.430 4.000 1619.470 4.280 ;
        RECT 1620.310 4.000 1635.570 4.280 ;
        RECT 1636.410 4.000 1648.450 4.280 ;
        RECT 1649.290 4.000 1661.330 4.280 ;
        RECT 1662.170 4.000 1674.210 4.280 ;
        RECT 1675.050 4.000 1690.310 4.280 ;
        RECT 1691.150 4.000 1703.190 4.280 ;
        RECT 1704.030 4.000 1716.070 4.280 ;
        RECT 1716.910 4.000 1732.170 4.280 ;
        RECT 1733.010 4.000 1745.050 4.280 ;
        RECT 1745.890 4.000 1757.930 4.280 ;
        RECT 1758.770 4.000 1770.810 4.280 ;
        RECT 1771.650 4.000 1786.910 4.280 ;
        RECT 1787.750 4.000 1799.790 4.280 ;
        RECT 1800.630 4.000 1812.670 4.280 ;
        RECT 1813.510 4.000 1825.550 4.280 ;
        RECT 1826.390 4.000 1841.650 4.280 ;
        RECT 1842.490 4.000 1854.530 4.280 ;
        RECT 1855.370 4.000 1867.410 4.280 ;
        RECT 1868.250 4.000 1883.510 4.280 ;
        RECT 1884.350 4.000 1896.390 4.280 ;
      LAYER met3 ;
        RECT 4.400 2393.240 1896.000 2394.105 ;
        RECT 4.000 2391.240 1896.000 2393.240 ;
        RECT 4.000 2389.840 1895.600 2391.240 ;
        RECT 4.000 2381.040 1896.000 2389.840 ;
        RECT 4.400 2379.640 1896.000 2381.040 ;
        RECT 4.000 2377.640 1896.000 2379.640 ;
        RECT 4.000 2376.240 1895.600 2377.640 ;
        RECT 4.000 2367.440 1896.000 2376.240 ;
        RECT 4.400 2366.040 1896.000 2367.440 ;
        RECT 4.000 2364.040 1896.000 2366.040 ;
        RECT 4.000 2362.640 1895.600 2364.040 ;
        RECT 4.000 2350.440 1896.000 2362.640 ;
        RECT 4.400 2349.040 1895.600 2350.440 ;
        RECT 4.000 2336.840 1896.000 2349.040 ;
        RECT 4.400 2335.440 1896.000 2336.840 ;
        RECT 4.000 2333.440 1896.000 2335.440 ;
        RECT 4.000 2332.040 1895.600 2333.440 ;
        RECT 4.000 2323.240 1896.000 2332.040 ;
        RECT 4.400 2321.840 1896.000 2323.240 ;
        RECT 4.000 2319.840 1896.000 2321.840 ;
        RECT 4.000 2318.440 1895.600 2319.840 ;
        RECT 4.000 2306.240 1896.000 2318.440 ;
        RECT 4.400 2304.840 1895.600 2306.240 ;
        RECT 4.000 2292.640 1896.000 2304.840 ;
        RECT 4.400 2291.240 1896.000 2292.640 ;
        RECT 4.000 2289.240 1896.000 2291.240 ;
        RECT 4.000 2287.840 1895.600 2289.240 ;
        RECT 4.000 2279.040 1896.000 2287.840 ;
        RECT 4.400 2277.640 1896.000 2279.040 ;
        RECT 4.000 2275.640 1896.000 2277.640 ;
        RECT 4.000 2274.240 1895.600 2275.640 ;
        RECT 4.000 2265.440 1896.000 2274.240 ;
        RECT 4.400 2264.040 1896.000 2265.440 ;
        RECT 4.000 2262.040 1896.000 2264.040 ;
        RECT 4.000 2260.640 1895.600 2262.040 ;
        RECT 4.000 2248.440 1896.000 2260.640 ;
        RECT 4.400 2247.040 1895.600 2248.440 ;
        RECT 4.000 2234.840 1896.000 2247.040 ;
        RECT 4.400 2233.440 1896.000 2234.840 ;
        RECT 4.000 2231.440 1896.000 2233.440 ;
        RECT 4.000 2230.040 1895.600 2231.440 ;
        RECT 4.000 2221.240 1896.000 2230.040 ;
        RECT 4.400 2219.840 1896.000 2221.240 ;
        RECT 4.000 2217.840 1896.000 2219.840 ;
        RECT 4.000 2216.440 1895.600 2217.840 ;
        RECT 4.000 2207.640 1896.000 2216.440 ;
        RECT 4.400 2206.240 1896.000 2207.640 ;
        RECT 4.000 2204.240 1896.000 2206.240 ;
        RECT 4.000 2202.840 1895.600 2204.240 ;
        RECT 4.000 2190.640 1896.000 2202.840 ;
        RECT 4.400 2189.240 1895.600 2190.640 ;
        RECT 4.000 2177.040 1896.000 2189.240 ;
        RECT 4.400 2175.640 1896.000 2177.040 ;
        RECT 4.000 2173.640 1896.000 2175.640 ;
        RECT 4.000 2172.240 1895.600 2173.640 ;
        RECT 4.000 2163.440 1896.000 2172.240 ;
        RECT 4.400 2162.040 1896.000 2163.440 ;
        RECT 4.000 2160.040 1896.000 2162.040 ;
        RECT 4.000 2158.640 1895.600 2160.040 ;
        RECT 4.000 2146.440 1896.000 2158.640 ;
        RECT 4.400 2145.040 1895.600 2146.440 ;
        RECT 4.000 2132.840 1896.000 2145.040 ;
        RECT 4.400 2131.440 1895.600 2132.840 ;
        RECT 4.000 2119.240 1896.000 2131.440 ;
        RECT 4.400 2117.840 1896.000 2119.240 ;
        RECT 4.000 2115.840 1896.000 2117.840 ;
        RECT 4.000 2114.440 1895.600 2115.840 ;
        RECT 4.000 2105.640 1896.000 2114.440 ;
        RECT 4.400 2104.240 1896.000 2105.640 ;
        RECT 4.000 2102.240 1896.000 2104.240 ;
        RECT 4.000 2100.840 1895.600 2102.240 ;
        RECT 4.000 2088.640 1896.000 2100.840 ;
        RECT 4.400 2087.240 1895.600 2088.640 ;
        RECT 4.000 2075.040 1896.000 2087.240 ;
        RECT 4.400 2073.640 1896.000 2075.040 ;
        RECT 4.000 2071.640 1896.000 2073.640 ;
        RECT 4.000 2070.240 1895.600 2071.640 ;
        RECT 4.000 2061.440 1896.000 2070.240 ;
        RECT 4.400 2060.040 1896.000 2061.440 ;
        RECT 4.000 2058.040 1896.000 2060.040 ;
        RECT 4.000 2056.640 1895.600 2058.040 ;
        RECT 4.000 2047.840 1896.000 2056.640 ;
        RECT 4.400 2046.440 1896.000 2047.840 ;
        RECT 4.000 2044.440 1896.000 2046.440 ;
        RECT 4.000 2043.040 1895.600 2044.440 ;
        RECT 4.000 2030.840 1896.000 2043.040 ;
        RECT 4.400 2029.440 1895.600 2030.840 ;
        RECT 4.000 2017.240 1896.000 2029.440 ;
        RECT 4.400 2015.840 1896.000 2017.240 ;
        RECT 4.000 2013.840 1896.000 2015.840 ;
        RECT 4.000 2012.440 1895.600 2013.840 ;
        RECT 4.000 2003.640 1896.000 2012.440 ;
        RECT 4.400 2002.240 1896.000 2003.640 ;
        RECT 4.000 2000.240 1896.000 2002.240 ;
        RECT 4.000 1998.840 1895.600 2000.240 ;
        RECT 4.000 1990.040 1896.000 1998.840 ;
        RECT 4.400 1988.640 1896.000 1990.040 ;
        RECT 4.000 1986.640 1896.000 1988.640 ;
        RECT 4.000 1985.240 1895.600 1986.640 ;
        RECT 4.000 1973.040 1896.000 1985.240 ;
        RECT 4.400 1971.640 1895.600 1973.040 ;
        RECT 4.000 1959.440 1896.000 1971.640 ;
        RECT 4.400 1958.040 1896.000 1959.440 ;
        RECT 4.000 1956.040 1896.000 1958.040 ;
        RECT 4.000 1954.640 1895.600 1956.040 ;
        RECT 4.000 1945.840 1896.000 1954.640 ;
        RECT 4.400 1944.440 1896.000 1945.840 ;
        RECT 4.000 1942.440 1896.000 1944.440 ;
        RECT 4.000 1941.040 1895.600 1942.440 ;
        RECT 4.000 1928.840 1896.000 1941.040 ;
        RECT 4.400 1927.440 1895.600 1928.840 ;
        RECT 4.000 1915.240 1896.000 1927.440 ;
        RECT 4.400 1913.840 1896.000 1915.240 ;
        RECT 4.000 1911.840 1896.000 1913.840 ;
        RECT 4.000 1910.440 1895.600 1911.840 ;
        RECT 4.000 1901.640 1896.000 1910.440 ;
        RECT 4.400 1900.240 1896.000 1901.640 ;
        RECT 4.000 1898.240 1896.000 1900.240 ;
        RECT 4.000 1896.840 1895.600 1898.240 ;
        RECT 4.000 1888.040 1896.000 1896.840 ;
        RECT 4.400 1886.640 1896.000 1888.040 ;
        RECT 4.000 1884.640 1896.000 1886.640 ;
        RECT 4.000 1883.240 1895.600 1884.640 ;
        RECT 4.000 1871.040 1896.000 1883.240 ;
        RECT 4.400 1869.640 1895.600 1871.040 ;
        RECT 4.000 1857.440 1896.000 1869.640 ;
        RECT 4.400 1856.040 1896.000 1857.440 ;
        RECT 4.000 1854.040 1896.000 1856.040 ;
        RECT 4.000 1852.640 1895.600 1854.040 ;
        RECT 4.000 1843.840 1896.000 1852.640 ;
        RECT 4.400 1842.440 1896.000 1843.840 ;
        RECT 4.000 1840.440 1896.000 1842.440 ;
        RECT 4.000 1839.040 1895.600 1840.440 ;
        RECT 4.000 1830.240 1896.000 1839.040 ;
        RECT 4.400 1828.840 1896.000 1830.240 ;
        RECT 4.000 1826.840 1896.000 1828.840 ;
        RECT 4.000 1825.440 1895.600 1826.840 ;
        RECT 4.000 1813.240 1896.000 1825.440 ;
        RECT 4.400 1811.840 1895.600 1813.240 ;
        RECT 4.000 1799.640 1896.000 1811.840 ;
        RECT 4.400 1798.240 1896.000 1799.640 ;
        RECT 4.000 1796.240 1896.000 1798.240 ;
        RECT 4.000 1794.840 1895.600 1796.240 ;
        RECT 4.000 1786.040 1896.000 1794.840 ;
        RECT 4.400 1784.640 1896.000 1786.040 ;
        RECT 4.000 1782.640 1896.000 1784.640 ;
        RECT 4.000 1781.240 1895.600 1782.640 ;
        RECT 4.000 1769.040 1896.000 1781.240 ;
        RECT 4.400 1767.640 1895.600 1769.040 ;
        RECT 4.000 1755.440 1896.000 1767.640 ;
        RECT 4.400 1754.040 1896.000 1755.440 ;
        RECT 4.000 1752.040 1896.000 1754.040 ;
        RECT 4.000 1750.640 1895.600 1752.040 ;
        RECT 4.000 1741.840 1896.000 1750.640 ;
        RECT 4.400 1740.440 1896.000 1741.840 ;
        RECT 4.000 1738.440 1896.000 1740.440 ;
        RECT 4.000 1737.040 1895.600 1738.440 ;
        RECT 4.000 1728.240 1896.000 1737.040 ;
        RECT 4.400 1726.840 1896.000 1728.240 ;
        RECT 4.000 1724.840 1896.000 1726.840 ;
        RECT 4.000 1723.440 1895.600 1724.840 ;
        RECT 4.000 1711.240 1896.000 1723.440 ;
        RECT 4.400 1709.840 1895.600 1711.240 ;
        RECT 4.000 1697.640 1896.000 1709.840 ;
        RECT 4.400 1696.240 1896.000 1697.640 ;
        RECT 4.000 1694.240 1896.000 1696.240 ;
        RECT 4.000 1692.840 1895.600 1694.240 ;
        RECT 4.000 1684.040 1896.000 1692.840 ;
        RECT 4.400 1682.640 1896.000 1684.040 ;
        RECT 4.000 1680.640 1896.000 1682.640 ;
        RECT 4.000 1679.240 1895.600 1680.640 ;
        RECT 4.000 1670.440 1896.000 1679.240 ;
        RECT 4.400 1669.040 1896.000 1670.440 ;
        RECT 4.000 1667.040 1896.000 1669.040 ;
        RECT 4.000 1665.640 1895.600 1667.040 ;
        RECT 4.000 1653.440 1896.000 1665.640 ;
        RECT 4.400 1652.040 1895.600 1653.440 ;
        RECT 4.000 1639.840 1896.000 1652.040 ;
        RECT 4.400 1638.440 1896.000 1639.840 ;
        RECT 4.000 1636.440 1896.000 1638.440 ;
        RECT 4.000 1635.040 1895.600 1636.440 ;
        RECT 4.000 1626.240 1896.000 1635.040 ;
        RECT 4.400 1624.840 1896.000 1626.240 ;
        RECT 4.000 1622.840 1896.000 1624.840 ;
        RECT 4.000 1621.440 1895.600 1622.840 ;
        RECT 4.000 1609.240 1896.000 1621.440 ;
        RECT 4.400 1607.840 1895.600 1609.240 ;
        RECT 4.000 1595.640 1896.000 1607.840 ;
        RECT 4.400 1594.240 1895.600 1595.640 ;
        RECT 4.000 1582.040 1896.000 1594.240 ;
        RECT 4.400 1580.640 1896.000 1582.040 ;
        RECT 4.000 1578.640 1896.000 1580.640 ;
        RECT 4.000 1577.240 1895.600 1578.640 ;
        RECT 4.000 1568.440 1896.000 1577.240 ;
        RECT 4.400 1567.040 1896.000 1568.440 ;
        RECT 4.000 1565.040 1896.000 1567.040 ;
        RECT 4.000 1563.640 1895.600 1565.040 ;
        RECT 4.000 1551.440 1896.000 1563.640 ;
        RECT 4.400 1550.040 1895.600 1551.440 ;
        RECT 4.000 1537.840 1896.000 1550.040 ;
        RECT 4.400 1536.440 1896.000 1537.840 ;
        RECT 4.000 1534.440 1896.000 1536.440 ;
        RECT 4.000 1533.040 1895.600 1534.440 ;
        RECT 4.000 1524.240 1896.000 1533.040 ;
        RECT 4.400 1522.840 1896.000 1524.240 ;
        RECT 4.000 1520.840 1896.000 1522.840 ;
        RECT 4.000 1519.440 1895.600 1520.840 ;
        RECT 4.000 1510.640 1896.000 1519.440 ;
        RECT 4.400 1509.240 1896.000 1510.640 ;
        RECT 4.000 1507.240 1896.000 1509.240 ;
        RECT 4.000 1505.840 1895.600 1507.240 ;
        RECT 4.000 1493.640 1896.000 1505.840 ;
        RECT 4.400 1492.240 1895.600 1493.640 ;
        RECT 4.000 1480.040 1896.000 1492.240 ;
        RECT 4.400 1478.640 1896.000 1480.040 ;
        RECT 4.000 1476.640 1896.000 1478.640 ;
        RECT 4.000 1475.240 1895.600 1476.640 ;
        RECT 4.000 1466.440 1896.000 1475.240 ;
        RECT 4.400 1465.040 1896.000 1466.440 ;
        RECT 4.000 1463.040 1896.000 1465.040 ;
        RECT 4.000 1461.640 1895.600 1463.040 ;
        RECT 4.000 1452.840 1896.000 1461.640 ;
        RECT 4.400 1451.440 1896.000 1452.840 ;
        RECT 4.000 1449.440 1896.000 1451.440 ;
        RECT 4.000 1448.040 1895.600 1449.440 ;
        RECT 4.000 1435.840 1896.000 1448.040 ;
        RECT 4.400 1434.440 1895.600 1435.840 ;
        RECT 4.000 1422.240 1896.000 1434.440 ;
        RECT 4.400 1420.840 1896.000 1422.240 ;
        RECT 4.000 1418.840 1896.000 1420.840 ;
        RECT 4.000 1417.440 1895.600 1418.840 ;
        RECT 4.000 1408.640 1896.000 1417.440 ;
        RECT 4.400 1407.240 1896.000 1408.640 ;
        RECT 4.000 1405.240 1896.000 1407.240 ;
        RECT 4.000 1403.840 1895.600 1405.240 ;
        RECT 4.000 1391.640 1896.000 1403.840 ;
        RECT 4.400 1390.240 1895.600 1391.640 ;
        RECT 4.000 1378.040 1896.000 1390.240 ;
        RECT 4.400 1376.640 1896.000 1378.040 ;
        RECT 4.000 1374.640 1896.000 1376.640 ;
        RECT 4.000 1373.240 1895.600 1374.640 ;
        RECT 4.000 1364.440 1896.000 1373.240 ;
        RECT 4.400 1363.040 1896.000 1364.440 ;
        RECT 4.000 1361.040 1896.000 1363.040 ;
        RECT 4.000 1359.640 1895.600 1361.040 ;
        RECT 4.000 1350.840 1896.000 1359.640 ;
        RECT 4.400 1349.440 1896.000 1350.840 ;
        RECT 4.000 1347.440 1896.000 1349.440 ;
        RECT 4.000 1346.040 1895.600 1347.440 ;
        RECT 4.000 1333.840 1896.000 1346.040 ;
        RECT 4.400 1332.440 1895.600 1333.840 ;
        RECT 4.000 1320.240 1896.000 1332.440 ;
        RECT 4.400 1318.840 1896.000 1320.240 ;
        RECT 4.000 1316.840 1896.000 1318.840 ;
        RECT 4.000 1315.440 1895.600 1316.840 ;
        RECT 4.000 1306.640 1896.000 1315.440 ;
        RECT 4.400 1305.240 1896.000 1306.640 ;
        RECT 4.000 1303.240 1896.000 1305.240 ;
        RECT 4.000 1301.840 1895.600 1303.240 ;
        RECT 4.000 1293.040 1896.000 1301.840 ;
        RECT 4.400 1291.640 1896.000 1293.040 ;
        RECT 4.000 1289.640 1896.000 1291.640 ;
        RECT 4.000 1288.240 1895.600 1289.640 ;
        RECT 4.000 1276.040 1896.000 1288.240 ;
        RECT 4.400 1274.640 1895.600 1276.040 ;
        RECT 4.000 1262.440 1896.000 1274.640 ;
        RECT 4.400 1261.040 1896.000 1262.440 ;
        RECT 4.000 1259.040 1896.000 1261.040 ;
        RECT 4.000 1257.640 1895.600 1259.040 ;
        RECT 4.000 1248.840 1896.000 1257.640 ;
        RECT 4.400 1247.440 1896.000 1248.840 ;
        RECT 4.000 1245.440 1896.000 1247.440 ;
        RECT 4.000 1244.040 1895.600 1245.440 ;
        RECT 4.000 1231.840 1896.000 1244.040 ;
        RECT 4.400 1230.440 1895.600 1231.840 ;
        RECT 4.000 1218.240 1896.000 1230.440 ;
        RECT 4.400 1216.840 1896.000 1218.240 ;
        RECT 4.000 1214.840 1896.000 1216.840 ;
        RECT 4.000 1213.440 1895.600 1214.840 ;
        RECT 4.000 1204.640 1896.000 1213.440 ;
        RECT 4.400 1203.240 1896.000 1204.640 ;
        RECT 4.000 1201.240 1896.000 1203.240 ;
        RECT 4.000 1199.840 1895.600 1201.240 ;
        RECT 4.000 1191.040 1896.000 1199.840 ;
        RECT 4.400 1189.640 1896.000 1191.040 ;
        RECT 4.000 1187.640 1896.000 1189.640 ;
        RECT 4.000 1186.240 1895.600 1187.640 ;
        RECT 4.000 1174.040 1896.000 1186.240 ;
        RECT 4.400 1172.640 1895.600 1174.040 ;
        RECT 4.000 1160.440 1896.000 1172.640 ;
        RECT 4.400 1159.040 1896.000 1160.440 ;
        RECT 4.000 1157.040 1896.000 1159.040 ;
        RECT 4.000 1155.640 1895.600 1157.040 ;
        RECT 4.000 1146.840 1896.000 1155.640 ;
        RECT 4.400 1145.440 1896.000 1146.840 ;
        RECT 4.000 1143.440 1896.000 1145.440 ;
        RECT 4.000 1142.040 1895.600 1143.440 ;
        RECT 4.000 1133.240 1896.000 1142.040 ;
        RECT 4.400 1131.840 1896.000 1133.240 ;
        RECT 4.000 1129.840 1896.000 1131.840 ;
        RECT 4.000 1128.440 1895.600 1129.840 ;
        RECT 4.000 1116.240 1896.000 1128.440 ;
        RECT 4.400 1114.840 1895.600 1116.240 ;
        RECT 4.000 1102.640 1896.000 1114.840 ;
        RECT 4.400 1101.240 1896.000 1102.640 ;
        RECT 4.000 1099.240 1896.000 1101.240 ;
        RECT 4.000 1097.840 1895.600 1099.240 ;
        RECT 4.000 1089.040 1896.000 1097.840 ;
        RECT 4.400 1087.640 1896.000 1089.040 ;
        RECT 4.000 1085.640 1896.000 1087.640 ;
        RECT 4.000 1084.240 1895.600 1085.640 ;
        RECT 4.000 1072.040 1896.000 1084.240 ;
        RECT 4.400 1070.640 1895.600 1072.040 ;
        RECT 4.000 1058.440 1896.000 1070.640 ;
        RECT 4.400 1057.040 1895.600 1058.440 ;
        RECT 4.000 1044.840 1896.000 1057.040 ;
        RECT 4.400 1043.440 1896.000 1044.840 ;
        RECT 4.000 1041.440 1896.000 1043.440 ;
        RECT 4.000 1040.040 1895.600 1041.440 ;
        RECT 4.000 1031.240 1896.000 1040.040 ;
        RECT 4.400 1029.840 1896.000 1031.240 ;
        RECT 4.000 1027.840 1896.000 1029.840 ;
        RECT 4.000 1026.440 1895.600 1027.840 ;
        RECT 4.000 1014.240 1896.000 1026.440 ;
        RECT 4.400 1012.840 1895.600 1014.240 ;
        RECT 4.000 1000.640 1896.000 1012.840 ;
        RECT 4.400 999.240 1896.000 1000.640 ;
        RECT 4.000 997.240 1896.000 999.240 ;
        RECT 4.000 995.840 1895.600 997.240 ;
        RECT 4.000 987.040 1896.000 995.840 ;
        RECT 4.400 985.640 1896.000 987.040 ;
        RECT 4.000 983.640 1896.000 985.640 ;
        RECT 4.000 982.240 1895.600 983.640 ;
        RECT 4.000 973.440 1896.000 982.240 ;
        RECT 4.400 972.040 1896.000 973.440 ;
        RECT 4.000 970.040 1896.000 972.040 ;
        RECT 4.000 968.640 1895.600 970.040 ;
        RECT 4.000 956.440 1896.000 968.640 ;
        RECT 4.400 955.040 1895.600 956.440 ;
        RECT 4.000 942.840 1896.000 955.040 ;
        RECT 4.400 941.440 1896.000 942.840 ;
        RECT 4.000 939.440 1896.000 941.440 ;
        RECT 4.000 938.040 1895.600 939.440 ;
        RECT 4.000 929.240 1896.000 938.040 ;
        RECT 4.400 927.840 1896.000 929.240 ;
        RECT 4.000 925.840 1896.000 927.840 ;
        RECT 4.000 924.440 1895.600 925.840 ;
        RECT 4.000 915.640 1896.000 924.440 ;
        RECT 4.400 914.240 1896.000 915.640 ;
        RECT 4.000 912.240 1896.000 914.240 ;
        RECT 4.000 910.840 1895.600 912.240 ;
        RECT 4.000 898.640 1896.000 910.840 ;
        RECT 4.400 897.240 1895.600 898.640 ;
        RECT 4.000 885.040 1896.000 897.240 ;
        RECT 4.400 883.640 1896.000 885.040 ;
        RECT 4.000 881.640 1896.000 883.640 ;
        RECT 4.000 880.240 1895.600 881.640 ;
        RECT 4.000 871.440 1896.000 880.240 ;
        RECT 4.400 870.040 1896.000 871.440 ;
        RECT 4.000 868.040 1896.000 870.040 ;
        RECT 4.000 866.640 1895.600 868.040 ;
        RECT 4.000 854.440 1896.000 866.640 ;
        RECT 4.400 853.040 1895.600 854.440 ;
        RECT 4.000 840.840 1896.000 853.040 ;
        RECT 4.400 839.440 1896.000 840.840 ;
        RECT 4.000 837.440 1896.000 839.440 ;
        RECT 4.000 836.040 1895.600 837.440 ;
        RECT 4.000 827.240 1896.000 836.040 ;
        RECT 4.400 825.840 1896.000 827.240 ;
        RECT 4.000 823.840 1896.000 825.840 ;
        RECT 4.000 822.440 1895.600 823.840 ;
        RECT 4.000 813.640 1896.000 822.440 ;
        RECT 4.400 812.240 1896.000 813.640 ;
        RECT 4.000 810.240 1896.000 812.240 ;
        RECT 4.000 808.840 1895.600 810.240 ;
        RECT 4.000 796.640 1896.000 808.840 ;
        RECT 4.400 795.240 1895.600 796.640 ;
        RECT 4.000 783.040 1896.000 795.240 ;
        RECT 4.400 781.640 1896.000 783.040 ;
        RECT 4.000 779.640 1896.000 781.640 ;
        RECT 4.000 778.240 1895.600 779.640 ;
        RECT 4.000 769.440 1896.000 778.240 ;
        RECT 4.400 768.040 1896.000 769.440 ;
        RECT 4.000 766.040 1896.000 768.040 ;
        RECT 4.000 764.640 1895.600 766.040 ;
        RECT 4.000 755.840 1896.000 764.640 ;
        RECT 4.400 754.440 1896.000 755.840 ;
        RECT 4.000 752.440 1896.000 754.440 ;
        RECT 4.000 751.040 1895.600 752.440 ;
        RECT 4.000 738.840 1896.000 751.040 ;
        RECT 4.400 737.440 1895.600 738.840 ;
        RECT 4.000 725.240 1896.000 737.440 ;
        RECT 4.400 723.840 1896.000 725.240 ;
        RECT 4.000 721.840 1896.000 723.840 ;
        RECT 4.000 720.440 1895.600 721.840 ;
        RECT 4.000 711.640 1896.000 720.440 ;
        RECT 4.400 710.240 1896.000 711.640 ;
        RECT 4.000 708.240 1896.000 710.240 ;
        RECT 4.000 706.840 1895.600 708.240 ;
        RECT 4.000 694.640 1896.000 706.840 ;
        RECT 4.400 693.240 1895.600 694.640 ;
        RECT 4.000 681.040 1896.000 693.240 ;
        RECT 4.400 679.640 1896.000 681.040 ;
        RECT 4.000 677.640 1896.000 679.640 ;
        RECT 4.000 676.240 1895.600 677.640 ;
        RECT 4.000 667.440 1896.000 676.240 ;
        RECT 4.400 666.040 1896.000 667.440 ;
        RECT 4.000 664.040 1896.000 666.040 ;
        RECT 4.000 662.640 1895.600 664.040 ;
        RECT 4.000 653.840 1896.000 662.640 ;
        RECT 4.400 652.440 1896.000 653.840 ;
        RECT 4.000 650.440 1896.000 652.440 ;
        RECT 4.000 649.040 1895.600 650.440 ;
        RECT 4.000 636.840 1896.000 649.040 ;
        RECT 4.400 635.440 1895.600 636.840 ;
        RECT 4.000 623.240 1896.000 635.440 ;
        RECT 4.400 621.840 1896.000 623.240 ;
        RECT 4.000 619.840 1896.000 621.840 ;
        RECT 4.000 618.440 1895.600 619.840 ;
        RECT 4.000 609.640 1896.000 618.440 ;
        RECT 4.400 608.240 1896.000 609.640 ;
        RECT 4.000 606.240 1896.000 608.240 ;
        RECT 4.000 604.840 1895.600 606.240 ;
        RECT 4.000 596.040 1896.000 604.840 ;
        RECT 4.400 594.640 1896.000 596.040 ;
        RECT 4.000 592.640 1896.000 594.640 ;
        RECT 4.000 591.240 1895.600 592.640 ;
        RECT 4.000 579.040 1896.000 591.240 ;
        RECT 4.400 577.640 1895.600 579.040 ;
        RECT 4.000 565.440 1896.000 577.640 ;
        RECT 4.400 564.040 1896.000 565.440 ;
        RECT 4.000 562.040 1896.000 564.040 ;
        RECT 4.000 560.640 1895.600 562.040 ;
        RECT 4.000 551.840 1896.000 560.640 ;
        RECT 4.400 550.440 1896.000 551.840 ;
        RECT 4.000 548.440 1896.000 550.440 ;
        RECT 4.000 547.040 1895.600 548.440 ;
        RECT 4.000 534.840 1896.000 547.040 ;
        RECT 4.400 533.440 1895.600 534.840 ;
        RECT 4.000 521.240 1896.000 533.440 ;
        RECT 4.400 519.840 1895.600 521.240 ;
        RECT 4.000 507.640 1896.000 519.840 ;
        RECT 4.400 506.240 1896.000 507.640 ;
        RECT 4.000 504.240 1896.000 506.240 ;
        RECT 4.000 502.840 1895.600 504.240 ;
        RECT 4.000 494.040 1896.000 502.840 ;
        RECT 4.400 492.640 1896.000 494.040 ;
        RECT 4.000 490.640 1896.000 492.640 ;
        RECT 4.000 489.240 1895.600 490.640 ;
        RECT 4.000 477.040 1896.000 489.240 ;
        RECT 4.400 475.640 1895.600 477.040 ;
        RECT 4.000 463.440 1896.000 475.640 ;
        RECT 4.400 462.040 1896.000 463.440 ;
        RECT 4.000 460.040 1896.000 462.040 ;
        RECT 4.000 458.640 1895.600 460.040 ;
        RECT 4.000 449.840 1896.000 458.640 ;
        RECT 4.400 448.440 1896.000 449.840 ;
        RECT 4.000 446.440 1896.000 448.440 ;
        RECT 4.000 445.040 1895.600 446.440 ;
        RECT 4.000 436.240 1896.000 445.040 ;
        RECT 4.400 434.840 1896.000 436.240 ;
        RECT 4.000 432.840 1896.000 434.840 ;
        RECT 4.000 431.440 1895.600 432.840 ;
        RECT 4.000 419.240 1896.000 431.440 ;
        RECT 4.400 417.840 1895.600 419.240 ;
        RECT 4.000 405.640 1896.000 417.840 ;
        RECT 4.400 404.240 1896.000 405.640 ;
        RECT 4.000 402.240 1896.000 404.240 ;
        RECT 4.000 400.840 1895.600 402.240 ;
        RECT 4.000 392.040 1896.000 400.840 ;
        RECT 4.400 390.640 1896.000 392.040 ;
        RECT 4.000 388.640 1896.000 390.640 ;
        RECT 4.000 387.240 1895.600 388.640 ;
        RECT 4.000 378.440 1896.000 387.240 ;
        RECT 4.400 377.040 1896.000 378.440 ;
        RECT 4.000 375.040 1896.000 377.040 ;
        RECT 4.000 373.640 1895.600 375.040 ;
        RECT 4.000 361.440 1896.000 373.640 ;
        RECT 4.400 360.040 1895.600 361.440 ;
        RECT 4.000 347.840 1896.000 360.040 ;
        RECT 4.400 346.440 1896.000 347.840 ;
        RECT 4.000 344.440 1896.000 346.440 ;
        RECT 4.000 343.040 1895.600 344.440 ;
        RECT 4.000 334.240 1896.000 343.040 ;
        RECT 4.400 332.840 1896.000 334.240 ;
        RECT 4.000 330.840 1896.000 332.840 ;
        RECT 4.000 329.440 1895.600 330.840 ;
        RECT 4.000 317.240 1896.000 329.440 ;
        RECT 4.400 315.840 1895.600 317.240 ;
        RECT 4.000 303.640 1896.000 315.840 ;
        RECT 4.400 302.240 1896.000 303.640 ;
        RECT 4.000 300.240 1896.000 302.240 ;
        RECT 4.000 298.840 1895.600 300.240 ;
        RECT 4.000 290.040 1896.000 298.840 ;
        RECT 4.400 288.640 1896.000 290.040 ;
        RECT 4.000 286.640 1896.000 288.640 ;
        RECT 4.000 285.240 1895.600 286.640 ;
        RECT 4.000 276.440 1896.000 285.240 ;
        RECT 4.400 275.040 1896.000 276.440 ;
        RECT 4.000 273.040 1896.000 275.040 ;
        RECT 4.000 271.640 1895.600 273.040 ;
        RECT 4.000 259.440 1896.000 271.640 ;
        RECT 4.400 258.040 1895.600 259.440 ;
        RECT 4.000 245.840 1896.000 258.040 ;
        RECT 4.400 244.440 1896.000 245.840 ;
        RECT 4.000 242.440 1896.000 244.440 ;
        RECT 4.000 241.040 1895.600 242.440 ;
        RECT 4.000 232.240 1896.000 241.040 ;
        RECT 4.400 230.840 1896.000 232.240 ;
        RECT 4.000 228.840 1896.000 230.840 ;
        RECT 4.000 227.440 1895.600 228.840 ;
        RECT 4.000 218.640 1896.000 227.440 ;
        RECT 4.400 217.240 1896.000 218.640 ;
        RECT 4.000 215.240 1896.000 217.240 ;
        RECT 4.000 213.840 1895.600 215.240 ;
        RECT 4.000 201.640 1896.000 213.840 ;
        RECT 4.400 200.240 1895.600 201.640 ;
        RECT 4.000 188.040 1896.000 200.240 ;
        RECT 4.400 186.640 1896.000 188.040 ;
        RECT 4.000 184.640 1896.000 186.640 ;
        RECT 4.000 183.240 1895.600 184.640 ;
        RECT 4.000 174.440 1896.000 183.240 ;
        RECT 4.400 173.040 1896.000 174.440 ;
        RECT 4.000 171.040 1896.000 173.040 ;
        RECT 4.000 169.640 1895.600 171.040 ;
        RECT 4.000 157.440 1896.000 169.640 ;
        RECT 4.400 156.040 1895.600 157.440 ;
        RECT 4.000 143.840 1896.000 156.040 ;
        RECT 4.400 142.440 1896.000 143.840 ;
        RECT 4.000 140.440 1896.000 142.440 ;
        RECT 4.000 139.040 1895.600 140.440 ;
        RECT 4.000 130.240 1896.000 139.040 ;
        RECT 4.400 128.840 1896.000 130.240 ;
        RECT 4.000 126.840 1896.000 128.840 ;
        RECT 4.000 125.440 1895.600 126.840 ;
        RECT 4.000 116.640 1896.000 125.440 ;
        RECT 4.400 115.240 1896.000 116.640 ;
        RECT 4.000 113.240 1896.000 115.240 ;
        RECT 4.000 111.840 1895.600 113.240 ;
        RECT 4.000 99.640 1896.000 111.840 ;
        RECT 4.400 98.240 1895.600 99.640 ;
        RECT 4.000 86.040 1896.000 98.240 ;
        RECT 4.400 84.640 1896.000 86.040 ;
        RECT 4.000 82.640 1896.000 84.640 ;
        RECT 4.000 81.240 1895.600 82.640 ;
        RECT 4.000 72.440 1896.000 81.240 ;
        RECT 4.400 71.040 1896.000 72.440 ;
        RECT 4.000 69.040 1896.000 71.040 ;
        RECT 4.000 67.640 1895.600 69.040 ;
        RECT 4.000 58.840 1896.000 67.640 ;
        RECT 4.400 57.440 1896.000 58.840 ;
        RECT 4.000 55.440 1896.000 57.440 ;
        RECT 4.000 54.040 1895.600 55.440 ;
        RECT 4.000 41.840 1896.000 54.040 ;
        RECT 4.400 40.440 1895.600 41.840 ;
        RECT 4.000 28.240 1896.000 40.440 ;
        RECT 4.400 26.840 1896.000 28.240 ;
        RECT 4.000 24.840 1896.000 26.840 ;
        RECT 4.000 23.440 1895.600 24.840 ;
        RECT 4.000 14.640 1896.000 23.440 ;
        RECT 4.400 13.240 1896.000 14.640 ;
        RECT 4.000 11.240 1896.000 13.240 ;
        RECT 4.000 10.375 1895.600 11.240 ;
      LAYER met4 ;
        RECT 1172.375 982.775 1172.640 994.665 ;
        RECT 1175.040 982.775 1175.465 994.665 ;
  END
END user_proj_systollic
END LIBRARY

